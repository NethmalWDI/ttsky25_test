magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -12993 -4583 -9047 1123
<< pwell >>
rect -126 234 586 326
rect -126 -2974 -34 234
rect 494 -2974 586 234
rect -126 -3106 586 -2974
<< psubdiff >>
rect -100 260 560 300
rect -100 -3000 -60 260
rect 520 -3000 560 260
rect -100 -3023 560 -3000
rect -100 -3057 -45 -3023
rect -11 -3057 23 -3023
rect 57 -3057 91 -3023
rect 125 -3057 159 -3023
rect 193 -3057 227 -3023
rect 261 -3057 295 -3023
rect 329 -3057 363 -3023
rect 397 -3057 431 -3023
rect 465 -3057 560 -3023
rect -100 -3080 560 -3057
<< nsubdiff >>
rect -12957 1053 -12873 1087
rect -12839 1053 -12805 1087
rect -12771 1053 -12737 1087
rect -12703 1053 -12669 1087
rect -12635 1053 -12601 1087
rect -12567 1053 -12533 1087
rect -12499 1053 -12465 1087
rect -12431 1053 -12397 1087
rect -12363 1053 -12329 1087
rect -12295 1053 -12261 1087
rect -12227 1053 -12193 1087
rect -12159 1053 -12125 1087
rect -12091 1053 -12057 1087
rect -12023 1053 -11989 1087
rect -11955 1053 -11921 1087
rect -11887 1053 -11853 1087
rect -11819 1053 -11785 1087
rect -11751 1053 -11717 1087
rect -11683 1053 -11649 1087
rect -11615 1053 -11581 1087
rect -11547 1053 -11513 1087
rect -11479 1053 -11445 1087
rect -11411 1053 -11377 1087
rect -11343 1053 -11309 1087
rect -11275 1053 -11241 1087
rect -11207 1053 -11173 1087
rect -11139 1053 -11105 1087
rect -11071 1053 -11037 1087
rect -11003 1053 -10969 1087
rect -10935 1053 -10901 1087
rect -10867 1053 -10833 1087
rect -10799 1053 -10765 1087
rect -10731 1053 -10697 1087
rect -10663 1053 -10629 1087
rect -10595 1053 -10561 1087
rect -10527 1053 -10493 1087
rect -10459 1053 -10425 1087
rect -10391 1053 -10357 1087
rect -10323 1053 -10289 1087
rect -10255 1053 -10221 1087
rect -10187 1053 -10153 1087
rect -10119 1053 -10085 1087
rect -10051 1053 -10017 1087
rect -9983 1053 -9949 1087
rect -9915 1053 -9881 1087
rect -9847 1053 -9813 1087
rect -9779 1053 -9745 1087
rect -9711 1053 -9677 1087
rect -9643 1053 -9609 1087
rect -9575 1053 -9541 1087
rect -9507 1053 -9473 1087
rect -9439 1053 -9405 1087
rect -9371 1053 -9337 1087
rect -9303 1053 -9269 1087
rect -9235 1053 -9201 1087
rect -9167 1053 -9083 1087
rect -12957 1007 -12923 1053
rect -12957 939 -12923 973
rect -12957 871 -12923 905
rect -12957 803 -12923 837
rect -12957 735 -12923 769
rect -12957 667 -12923 701
rect -12957 599 -12923 633
rect -12957 531 -12923 565
rect -12957 463 -12923 497
rect -12957 395 -12923 429
rect -12957 327 -12923 361
rect -12957 259 -12923 293
rect -12957 191 -12923 225
rect -12957 123 -12923 157
rect -12957 55 -12923 89
rect -12957 -13 -12923 21
rect -12957 -81 -12923 -47
rect -12957 -149 -12923 -115
rect -12957 -217 -12923 -183
rect -12957 -285 -12923 -251
rect -12957 -353 -12923 -319
rect -12957 -421 -12923 -387
rect -12957 -489 -12923 -455
rect -12957 -557 -12923 -523
rect -12957 -625 -12923 -591
rect -12957 -693 -12923 -659
rect -12957 -761 -12923 -727
rect -12957 -829 -12923 -795
rect -12957 -897 -12923 -863
rect -12957 -965 -12923 -931
rect -12957 -1033 -12923 -999
rect -12957 -1101 -12923 -1067
rect -12957 -1169 -12923 -1135
rect -12957 -1237 -12923 -1203
rect -12957 -1305 -12923 -1271
rect -12957 -1373 -12923 -1339
rect -12957 -1441 -12923 -1407
rect -12957 -1509 -12923 -1475
rect -12957 -1577 -12923 -1543
rect -12957 -1645 -12923 -1611
rect -12957 -1713 -12923 -1679
rect -12957 -1781 -12923 -1747
rect -12957 -1849 -12923 -1815
rect -12957 -1917 -12923 -1883
rect -12957 -1985 -12923 -1951
rect -12957 -2053 -12923 -2019
rect -12957 -2121 -12923 -2087
rect -12957 -2189 -12923 -2155
rect -12957 -2257 -12923 -2223
rect -12957 -2325 -12923 -2291
rect -12957 -2393 -12923 -2359
rect -12957 -2461 -12923 -2427
rect -12957 -2529 -12923 -2495
rect -12957 -2597 -12923 -2563
rect -12957 -2665 -12923 -2631
rect -12957 -2733 -12923 -2699
rect -12957 -2801 -12923 -2767
rect -12957 -2869 -12923 -2835
rect -12957 -2937 -12923 -2903
rect -12957 -3005 -12923 -2971
rect -12957 -3073 -12923 -3039
rect -12957 -3141 -12923 -3107
rect -12957 -3209 -12923 -3175
rect -12957 -3277 -12923 -3243
rect -12957 -3345 -12923 -3311
rect -12957 -3413 -12923 -3379
rect -12957 -3481 -12923 -3447
rect -12957 -3549 -12923 -3515
rect -12957 -3617 -12923 -3583
rect -12957 -3685 -12923 -3651
rect -12957 -3753 -12923 -3719
rect -12957 -3821 -12923 -3787
rect -12957 -3889 -12923 -3855
rect -12957 -3957 -12923 -3923
rect -12957 -4025 -12923 -3991
rect -12957 -4093 -12923 -4059
rect -12957 -4161 -12923 -4127
rect -12957 -4229 -12923 -4195
rect -12957 -4297 -12923 -4263
rect -12957 -4365 -12923 -4331
rect -12957 -4433 -12923 -4399
rect -12957 -4513 -12923 -4467
rect -9117 1007 -9083 1053
rect -9117 939 -9083 973
rect -9117 871 -9083 905
rect -9117 803 -9083 837
rect -9117 735 -9083 769
rect -9117 667 -9083 701
rect -9117 599 -9083 633
rect -9117 531 -9083 565
rect -9117 463 -9083 497
rect -9117 395 -9083 429
rect -9117 327 -9083 361
rect -9117 259 -9083 293
rect -9117 191 -9083 225
rect -9117 123 -9083 157
rect -9117 55 -9083 89
rect -9117 -13 -9083 21
rect -9117 -81 -9083 -47
rect -9117 -149 -9083 -115
rect -9117 -217 -9083 -183
rect -9117 -285 -9083 -251
rect -9117 -353 -9083 -319
rect -9117 -421 -9083 -387
rect -9117 -489 -9083 -455
rect -9117 -557 -9083 -523
rect -9117 -625 -9083 -591
rect -9117 -693 -9083 -659
rect -9117 -761 -9083 -727
rect -9117 -829 -9083 -795
rect -9117 -897 -9083 -863
rect -9117 -965 -9083 -931
rect -9117 -1033 -9083 -999
rect -9117 -1101 -9083 -1067
rect -9117 -1169 -9083 -1135
rect -9117 -1237 -9083 -1203
rect -9117 -1305 -9083 -1271
rect -9117 -1373 -9083 -1339
rect -9117 -1441 -9083 -1407
rect -9117 -1509 -9083 -1475
rect -9117 -1577 -9083 -1543
rect -9117 -1645 -9083 -1611
rect -9117 -1713 -9083 -1679
rect -9117 -1781 -9083 -1747
rect -9117 -1849 -9083 -1815
rect -9117 -1917 -9083 -1883
rect -9117 -1985 -9083 -1951
rect -9117 -2053 -9083 -2019
rect -9117 -2121 -9083 -2087
rect -9117 -2189 -9083 -2155
rect -9117 -2257 -9083 -2223
rect -9117 -2325 -9083 -2291
rect -9117 -2393 -9083 -2359
rect -9117 -2461 -9083 -2427
rect -9117 -2529 -9083 -2495
rect -9117 -2597 -9083 -2563
rect -9117 -2665 -9083 -2631
rect -9117 -2733 -9083 -2699
rect -9117 -2801 -9083 -2767
rect -9117 -2869 -9083 -2835
rect -9117 -2937 -9083 -2903
rect -9117 -3005 -9083 -2971
rect -9117 -3073 -9083 -3039
rect -9117 -3141 -9083 -3107
rect -9117 -3209 -9083 -3175
rect -9117 -3277 -9083 -3243
rect -9117 -3345 -9083 -3311
rect -9117 -3413 -9083 -3379
rect -9117 -3481 -9083 -3447
rect -9117 -3549 -9083 -3515
rect -9117 -3617 -9083 -3583
rect -9117 -3685 -9083 -3651
rect -9117 -3753 -9083 -3719
rect -9117 -3821 -9083 -3787
rect -9117 -3889 -9083 -3855
rect -9117 -3957 -9083 -3923
rect -9117 -4025 -9083 -3991
rect -9117 -4093 -9083 -4059
rect -9117 -4161 -9083 -4127
rect -9117 -4229 -9083 -4195
rect -9117 -4297 -9083 -4263
rect -9117 -4365 -9083 -4331
rect -9117 -4433 -9083 -4399
rect -9117 -4513 -9083 -4467
rect -12957 -4547 -12873 -4513
rect -12839 -4547 -12805 -4513
rect -12771 -4547 -12737 -4513
rect -12703 -4547 -12669 -4513
rect -12635 -4547 -12601 -4513
rect -12567 -4547 -12533 -4513
rect -12499 -4547 -12465 -4513
rect -12431 -4547 -12397 -4513
rect -12363 -4547 -12329 -4513
rect -12295 -4547 -12261 -4513
rect -12227 -4547 -12193 -4513
rect -12159 -4547 -12125 -4513
rect -12091 -4547 -12057 -4513
rect -12023 -4547 -11989 -4513
rect -11955 -4547 -11921 -4513
rect -11887 -4547 -11853 -4513
rect -11819 -4547 -11785 -4513
rect -11751 -4547 -11717 -4513
rect -11683 -4547 -11649 -4513
rect -11615 -4547 -11581 -4513
rect -11547 -4547 -11513 -4513
rect -11479 -4547 -11445 -4513
rect -11411 -4547 -11377 -4513
rect -11343 -4547 -11309 -4513
rect -11275 -4547 -11241 -4513
rect -11207 -4547 -11173 -4513
rect -11139 -4547 -11105 -4513
rect -11071 -4547 -11037 -4513
rect -11003 -4547 -10969 -4513
rect -10935 -4547 -10901 -4513
rect -10867 -4547 -10833 -4513
rect -10799 -4547 -10765 -4513
rect -10731 -4547 -10697 -4513
rect -10663 -4547 -10629 -4513
rect -10595 -4547 -10561 -4513
rect -10527 -4547 -10493 -4513
rect -10459 -4547 -10425 -4513
rect -10391 -4547 -10357 -4513
rect -10323 -4547 -10289 -4513
rect -10255 -4547 -10221 -4513
rect -10187 -4547 -10153 -4513
rect -10119 -4547 -10085 -4513
rect -10051 -4547 -10017 -4513
rect -9983 -4547 -9949 -4513
rect -9915 -4547 -9881 -4513
rect -9847 -4547 -9813 -4513
rect -9779 -4547 -9745 -4513
rect -9711 -4547 -9677 -4513
rect -9643 -4547 -9609 -4513
rect -9575 -4547 -9541 -4513
rect -9507 -4547 -9473 -4513
rect -9439 -4547 -9405 -4513
rect -9371 -4547 -9337 -4513
rect -9303 -4547 -9269 -4513
rect -9235 -4547 -9201 -4513
rect -9167 -4547 -9083 -4513
<< psubdiffcont >>
rect -45 -3057 -11 -3023
rect 23 -3057 57 -3023
rect 91 -3057 125 -3023
rect 159 -3057 193 -3023
rect 227 -3057 261 -3023
rect 295 -3057 329 -3023
rect 363 -3057 397 -3023
rect 431 -3057 465 -3023
<< nsubdiffcont >>
rect -12873 1053 -12839 1087
rect -12805 1053 -12771 1087
rect -12737 1053 -12703 1087
rect -12669 1053 -12635 1087
rect -12601 1053 -12567 1087
rect -12533 1053 -12499 1087
rect -12465 1053 -12431 1087
rect -12397 1053 -12363 1087
rect -12329 1053 -12295 1087
rect -12261 1053 -12227 1087
rect -12193 1053 -12159 1087
rect -12125 1053 -12091 1087
rect -12057 1053 -12023 1087
rect -11989 1053 -11955 1087
rect -11921 1053 -11887 1087
rect -11853 1053 -11819 1087
rect -11785 1053 -11751 1087
rect -11717 1053 -11683 1087
rect -11649 1053 -11615 1087
rect -11581 1053 -11547 1087
rect -11513 1053 -11479 1087
rect -11445 1053 -11411 1087
rect -11377 1053 -11343 1087
rect -11309 1053 -11275 1087
rect -11241 1053 -11207 1087
rect -11173 1053 -11139 1087
rect -11105 1053 -11071 1087
rect -11037 1053 -11003 1087
rect -10969 1053 -10935 1087
rect -10901 1053 -10867 1087
rect -10833 1053 -10799 1087
rect -10765 1053 -10731 1087
rect -10697 1053 -10663 1087
rect -10629 1053 -10595 1087
rect -10561 1053 -10527 1087
rect -10493 1053 -10459 1087
rect -10425 1053 -10391 1087
rect -10357 1053 -10323 1087
rect -10289 1053 -10255 1087
rect -10221 1053 -10187 1087
rect -10153 1053 -10119 1087
rect -10085 1053 -10051 1087
rect -10017 1053 -9983 1087
rect -9949 1053 -9915 1087
rect -9881 1053 -9847 1087
rect -9813 1053 -9779 1087
rect -9745 1053 -9711 1087
rect -9677 1053 -9643 1087
rect -9609 1053 -9575 1087
rect -9541 1053 -9507 1087
rect -9473 1053 -9439 1087
rect -9405 1053 -9371 1087
rect -9337 1053 -9303 1087
rect -9269 1053 -9235 1087
rect -9201 1053 -9167 1087
rect -12957 973 -12923 1007
rect -12957 905 -12923 939
rect -12957 837 -12923 871
rect -12957 769 -12923 803
rect -12957 701 -12923 735
rect -12957 633 -12923 667
rect -12957 565 -12923 599
rect -12957 497 -12923 531
rect -12957 429 -12923 463
rect -12957 361 -12923 395
rect -12957 293 -12923 327
rect -12957 225 -12923 259
rect -12957 157 -12923 191
rect -12957 89 -12923 123
rect -12957 21 -12923 55
rect -12957 -47 -12923 -13
rect -12957 -115 -12923 -81
rect -12957 -183 -12923 -149
rect -12957 -251 -12923 -217
rect -12957 -319 -12923 -285
rect -12957 -387 -12923 -353
rect -12957 -455 -12923 -421
rect -12957 -523 -12923 -489
rect -12957 -591 -12923 -557
rect -12957 -659 -12923 -625
rect -12957 -727 -12923 -693
rect -12957 -795 -12923 -761
rect -12957 -863 -12923 -829
rect -12957 -931 -12923 -897
rect -12957 -999 -12923 -965
rect -12957 -1067 -12923 -1033
rect -12957 -1135 -12923 -1101
rect -12957 -1203 -12923 -1169
rect -12957 -1271 -12923 -1237
rect -12957 -1339 -12923 -1305
rect -12957 -1407 -12923 -1373
rect -12957 -1475 -12923 -1441
rect -12957 -1543 -12923 -1509
rect -12957 -1611 -12923 -1577
rect -12957 -1679 -12923 -1645
rect -12957 -1747 -12923 -1713
rect -12957 -1815 -12923 -1781
rect -12957 -1883 -12923 -1849
rect -12957 -1951 -12923 -1917
rect -12957 -2019 -12923 -1985
rect -12957 -2087 -12923 -2053
rect -12957 -2155 -12923 -2121
rect -12957 -2223 -12923 -2189
rect -12957 -2291 -12923 -2257
rect -12957 -2359 -12923 -2325
rect -12957 -2427 -12923 -2393
rect -12957 -2495 -12923 -2461
rect -12957 -2563 -12923 -2529
rect -12957 -2631 -12923 -2597
rect -12957 -2699 -12923 -2665
rect -12957 -2767 -12923 -2733
rect -12957 -2835 -12923 -2801
rect -12957 -2903 -12923 -2869
rect -12957 -2971 -12923 -2937
rect -12957 -3039 -12923 -3005
rect -12957 -3107 -12923 -3073
rect -12957 -3175 -12923 -3141
rect -12957 -3243 -12923 -3209
rect -12957 -3311 -12923 -3277
rect -12957 -3379 -12923 -3345
rect -12957 -3447 -12923 -3413
rect -12957 -3515 -12923 -3481
rect -12957 -3583 -12923 -3549
rect -12957 -3651 -12923 -3617
rect -12957 -3719 -12923 -3685
rect -12957 -3787 -12923 -3753
rect -12957 -3855 -12923 -3821
rect -12957 -3923 -12923 -3889
rect -12957 -3991 -12923 -3957
rect -12957 -4059 -12923 -4025
rect -12957 -4127 -12923 -4093
rect -12957 -4195 -12923 -4161
rect -12957 -4263 -12923 -4229
rect -12957 -4331 -12923 -4297
rect -12957 -4399 -12923 -4365
rect -12957 -4467 -12923 -4433
rect -9117 973 -9083 1007
rect -9117 905 -9083 939
rect -9117 837 -9083 871
rect -9117 769 -9083 803
rect -9117 701 -9083 735
rect -9117 633 -9083 667
rect -9117 565 -9083 599
rect -9117 497 -9083 531
rect -9117 429 -9083 463
rect -9117 361 -9083 395
rect -9117 293 -9083 327
rect -9117 225 -9083 259
rect -9117 157 -9083 191
rect -9117 89 -9083 123
rect -9117 21 -9083 55
rect -9117 -47 -9083 -13
rect -9117 -115 -9083 -81
rect -9117 -183 -9083 -149
rect -9117 -251 -9083 -217
rect -9117 -319 -9083 -285
rect -9117 -387 -9083 -353
rect -9117 -455 -9083 -421
rect -9117 -523 -9083 -489
rect -9117 -591 -9083 -557
rect -9117 -659 -9083 -625
rect -9117 -727 -9083 -693
rect -9117 -795 -9083 -761
rect -9117 -863 -9083 -829
rect -9117 -931 -9083 -897
rect -9117 -999 -9083 -965
rect -9117 -1067 -9083 -1033
rect -9117 -1135 -9083 -1101
rect -9117 -1203 -9083 -1169
rect -9117 -1271 -9083 -1237
rect -9117 -1339 -9083 -1305
rect -9117 -1407 -9083 -1373
rect -9117 -1475 -9083 -1441
rect -9117 -1543 -9083 -1509
rect -9117 -1611 -9083 -1577
rect -9117 -1679 -9083 -1645
rect -9117 -1747 -9083 -1713
rect -9117 -1815 -9083 -1781
rect -9117 -1883 -9083 -1849
rect -9117 -1951 -9083 -1917
rect -9117 -2019 -9083 -1985
rect -9117 -2087 -9083 -2053
rect -9117 -2155 -9083 -2121
rect -9117 -2223 -9083 -2189
rect -9117 -2291 -9083 -2257
rect -9117 -2359 -9083 -2325
rect -9117 -2427 -9083 -2393
rect -9117 -2495 -9083 -2461
rect -9117 -2563 -9083 -2529
rect -9117 -2631 -9083 -2597
rect -9117 -2699 -9083 -2665
rect -9117 -2767 -9083 -2733
rect -9117 -2835 -9083 -2801
rect -9117 -2903 -9083 -2869
rect -9117 -2971 -9083 -2937
rect -9117 -3039 -9083 -3005
rect -9117 -3107 -9083 -3073
rect -9117 -3175 -9083 -3141
rect -9117 -3243 -9083 -3209
rect -9117 -3311 -9083 -3277
rect -9117 -3379 -9083 -3345
rect -9117 -3447 -9083 -3413
rect -9117 -3515 -9083 -3481
rect -9117 -3583 -9083 -3549
rect -9117 -3651 -9083 -3617
rect -9117 -3719 -9083 -3685
rect -9117 -3787 -9083 -3753
rect -9117 -3855 -9083 -3821
rect -9117 -3923 -9083 -3889
rect -9117 -3991 -9083 -3957
rect -9117 -4059 -9083 -4025
rect -9117 -4127 -9083 -4093
rect -9117 -4195 -9083 -4161
rect -9117 -4263 -9083 -4229
rect -9117 -4331 -9083 -4297
rect -9117 -4399 -9083 -4365
rect -9117 -4467 -9083 -4433
rect -12873 -4547 -12839 -4513
rect -12805 -4547 -12771 -4513
rect -12737 -4547 -12703 -4513
rect -12669 -4547 -12635 -4513
rect -12601 -4547 -12567 -4513
rect -12533 -4547 -12499 -4513
rect -12465 -4547 -12431 -4513
rect -12397 -4547 -12363 -4513
rect -12329 -4547 -12295 -4513
rect -12261 -4547 -12227 -4513
rect -12193 -4547 -12159 -4513
rect -12125 -4547 -12091 -4513
rect -12057 -4547 -12023 -4513
rect -11989 -4547 -11955 -4513
rect -11921 -4547 -11887 -4513
rect -11853 -4547 -11819 -4513
rect -11785 -4547 -11751 -4513
rect -11717 -4547 -11683 -4513
rect -11649 -4547 -11615 -4513
rect -11581 -4547 -11547 -4513
rect -11513 -4547 -11479 -4513
rect -11445 -4547 -11411 -4513
rect -11377 -4547 -11343 -4513
rect -11309 -4547 -11275 -4513
rect -11241 -4547 -11207 -4513
rect -11173 -4547 -11139 -4513
rect -11105 -4547 -11071 -4513
rect -11037 -4547 -11003 -4513
rect -10969 -4547 -10935 -4513
rect -10901 -4547 -10867 -4513
rect -10833 -4547 -10799 -4513
rect -10765 -4547 -10731 -4513
rect -10697 -4547 -10663 -4513
rect -10629 -4547 -10595 -4513
rect -10561 -4547 -10527 -4513
rect -10493 -4547 -10459 -4513
rect -10425 -4547 -10391 -4513
rect -10357 -4547 -10323 -4513
rect -10289 -4547 -10255 -4513
rect -10221 -4547 -10187 -4513
rect -10153 -4547 -10119 -4513
rect -10085 -4547 -10051 -4513
rect -10017 -4547 -9983 -4513
rect -9949 -4547 -9915 -4513
rect -9881 -4547 -9847 -4513
rect -9813 -4547 -9779 -4513
rect -9745 -4547 -9711 -4513
rect -9677 -4547 -9643 -4513
rect -9609 -4547 -9575 -4513
rect -9541 -4547 -9507 -4513
rect -9473 -4547 -9439 -4513
rect -9405 -4547 -9371 -4513
rect -9337 -4547 -9303 -4513
rect -9269 -4547 -9235 -4513
rect -9201 -4547 -9167 -4513
<< locali >>
rect -12957 1053 -12873 1087
rect -12839 1053 -12805 1087
rect -12771 1053 -12737 1087
rect -12703 1053 -12669 1087
rect -12635 1053 -12601 1087
rect -12567 1053 -12533 1087
rect -12499 1053 -12465 1087
rect -12431 1053 -12397 1087
rect -12363 1053 -12329 1087
rect -12295 1053 -12261 1087
rect -12227 1053 -12193 1087
rect -12159 1053 -12125 1087
rect -12091 1053 -12057 1087
rect -12023 1053 -11989 1087
rect -11955 1053 -11921 1087
rect -11887 1053 -11853 1087
rect -11819 1053 -11785 1087
rect -11751 1053 -11717 1087
rect -11683 1053 -11649 1087
rect -11615 1053 -11581 1087
rect -11547 1053 -11513 1087
rect -11479 1053 -11445 1087
rect -11411 1053 -11377 1087
rect -11343 1053 -11309 1087
rect -11275 1053 -11241 1087
rect -11207 1053 -11173 1087
rect -11139 1053 -11105 1087
rect -11071 1053 -11037 1087
rect -11003 1053 -10969 1087
rect -10935 1053 -10901 1087
rect -10867 1053 -10833 1087
rect -10799 1053 -10765 1087
rect -10731 1053 -10697 1087
rect -10663 1053 -10629 1087
rect -10595 1053 -10561 1087
rect -10527 1053 -10493 1087
rect -10459 1053 -10425 1087
rect -10391 1053 -10357 1087
rect -10323 1053 -10289 1087
rect -10255 1053 -10221 1087
rect -10187 1053 -10153 1087
rect -10119 1053 -10085 1087
rect -10051 1053 -10017 1087
rect -9983 1053 -9949 1087
rect -9915 1053 -9881 1087
rect -9847 1053 -9813 1087
rect -9779 1053 -9745 1087
rect -9711 1053 -9677 1087
rect -9643 1053 -9609 1087
rect -9575 1053 -9541 1087
rect -9507 1053 -9473 1087
rect -9439 1053 -9405 1087
rect -9371 1053 -9337 1087
rect -9303 1053 -9269 1087
rect -9235 1053 -9201 1087
rect -9167 1053 -9083 1087
rect -12957 1007 -12923 1053
rect -12957 939 -12923 973
rect -12957 871 -12923 905
rect -12957 803 -12923 837
rect -12957 735 -12923 769
rect -12957 667 -12923 701
rect -12957 599 -12923 633
rect -12957 531 -12923 565
rect -12957 463 -12923 497
rect -12957 395 -12923 429
rect -12957 327 -12923 361
rect -12957 259 -12923 293
rect -12957 191 -12923 225
rect -12957 123 -12923 157
rect -12957 55 -12923 89
rect -12957 -13 -12923 21
rect -12957 -81 -12923 -47
rect -12957 -149 -12923 -115
rect -12957 -217 -12923 -183
rect -12957 -285 -12923 -251
rect -12957 -353 -12923 -319
rect -12957 -421 -12923 -387
rect -12957 -489 -12923 -455
rect -12957 -557 -12923 -523
rect -12957 -625 -12923 -591
rect -12957 -693 -12923 -659
rect -12957 -761 -12923 -727
rect -12957 -829 -12923 -795
rect -12957 -897 -12923 -863
rect -12957 -965 -12923 -931
rect -12957 -1033 -12923 -999
rect -12957 -1101 -12923 -1067
rect -12957 -1169 -12923 -1135
rect -12957 -1237 -12923 -1203
rect -12957 -1305 -12923 -1271
rect -12957 -1373 -12923 -1339
rect -12957 -1441 -12923 -1407
rect -12957 -1509 -12923 -1475
rect -12957 -1577 -12923 -1543
rect -12957 -1645 -12923 -1611
rect -12957 -1713 -12923 -1679
rect -12957 -1781 -12923 -1747
rect -12957 -1849 -12923 -1815
rect -12957 -1917 -12923 -1883
rect -12957 -1985 -12923 -1951
rect -12957 -2053 -12923 -2019
rect -12957 -2121 -12923 -2087
rect -12957 -2189 -12923 -2155
rect -12957 -2257 -12923 -2223
rect -12957 -2325 -12923 -2291
rect -12957 -2393 -12923 -2359
rect -12957 -2461 -12923 -2427
rect -12957 -2529 -12923 -2495
rect -12957 -2597 -12923 -2563
rect -12957 -2665 -12923 -2631
rect -12957 -2733 -12923 -2699
rect -12957 -2801 -12923 -2767
rect -12957 -2869 -12923 -2835
rect -12957 -2937 -12923 -2903
rect -12957 -3005 -12923 -2971
rect -12957 -3073 -12923 -3039
rect -12957 -3141 -12923 -3107
rect -12957 -3209 -12923 -3175
rect -12957 -3277 -12923 -3243
rect -12957 -3345 -12923 -3311
rect -12957 -3413 -12923 -3379
rect -12957 -3481 -12923 -3447
rect -12957 -3549 -12923 -3515
rect -12957 -3617 -12923 -3583
rect -12957 -3685 -12923 -3651
rect -12957 -3753 -12923 -3719
rect -12957 -3821 -12923 -3787
rect -12957 -3889 -12923 -3855
rect -12957 -3957 -12923 -3923
rect -12957 -4025 -12923 -3991
rect -12957 -4093 -12923 -4059
rect -12957 -4161 -12923 -4127
rect -12957 -4229 -12923 -4195
rect -12957 -4297 -12923 -4263
rect -12957 -4365 -12923 -4331
rect -12957 -4433 -12923 -4399
rect -12957 -4513 -12923 -4467
rect -9117 1007 -9083 1053
rect -9117 939 -9083 973
rect -9117 871 -9083 905
rect -9117 803 -9083 837
rect -9117 735 -9083 769
rect -9117 667 -9083 701
rect -9117 599 -9083 633
rect -9117 531 -9083 565
rect -9117 463 -9083 497
rect -9117 395 -9083 429
rect -9117 327 -9083 361
rect -9117 259 -9083 293
rect -9117 191 -9083 225
rect -9117 123 -9083 157
rect -9117 55 -9083 89
rect -9117 -13 -9083 21
rect -9117 -81 -9083 -47
rect -9117 -149 -9083 -115
rect -9117 -217 -9083 -183
rect -9117 -285 -9083 -251
rect -9117 -353 -9083 -319
rect -9117 -421 -9083 -387
rect -9117 -489 -9083 -455
rect -9117 -557 -9083 -523
rect -9117 -625 -9083 -591
rect -9117 -693 -9083 -659
rect -9117 -761 -9083 -727
rect -9117 -829 -9083 -795
rect -9117 -897 -9083 -863
rect -9117 -965 -9083 -931
rect -9117 -1033 -9083 -999
rect -9117 -1101 -9083 -1067
rect -9117 -1169 -9083 -1135
rect -9117 -1237 -9083 -1203
rect -9117 -1305 -9083 -1271
rect -9117 -1373 -9083 -1339
rect -9117 -1441 -9083 -1407
rect -9117 -1509 -9083 -1475
rect -9117 -1577 -9083 -1543
rect -9117 -1645 -9083 -1611
rect -9117 -1713 -9083 -1679
rect -9117 -1781 -9083 -1747
rect -9117 -1849 -9083 -1815
rect -9117 -1917 -9083 -1883
rect -9117 -1985 -9083 -1951
rect -9117 -2053 -9083 -2019
rect -9117 -2121 -9083 -2087
rect -9117 -2189 -9083 -2155
rect -9117 -2257 -9083 -2223
rect -9117 -2325 -9083 -2291
rect -9117 -2393 -9083 -2359
rect -9117 -2461 -9083 -2427
rect -9117 -2529 -9083 -2495
rect -9117 -2597 -9083 -2563
rect -9117 -2665 -9083 -2631
rect -9117 -2733 -9083 -2699
rect -9117 -2801 -9083 -2767
rect -9117 -2869 -9083 -2835
rect -9117 -2937 -9083 -2903
rect -9117 -3005 -9083 -2971
rect -9117 -3073 -9083 -3039
rect -100 260 560 300
rect -100 -3000 -60 260
rect 520 -3000 560 260
rect -100 -3023 560 -3000
rect -100 -3057 -59 -3023
rect -11 -3057 13 -3023
rect 57 -3057 85 -3023
rect 125 -3057 157 -3023
rect 193 -3057 227 -3023
rect 263 -3057 295 -3023
rect 335 -3057 363 -3023
rect 407 -3057 431 -3023
rect 479 -3057 560 -3023
rect -100 -3080 560 -3057
rect -9117 -3141 -9083 -3107
rect -9117 -3209 -9083 -3175
rect -9117 -3277 -9083 -3243
rect -9117 -3345 -9083 -3311
rect -9117 -3413 -9083 -3379
rect -9117 -3481 -9083 -3447
rect -9117 -3549 -9083 -3515
rect -9117 -3617 -9083 -3583
rect -9117 -3685 -9083 -3651
rect -9117 -3753 -9083 -3719
rect -9117 -3821 -9083 -3787
rect -9117 -3889 -9083 -3855
rect -9117 -3957 -9083 -3923
rect -9117 -4025 -9083 -3991
rect -9117 -4093 -9083 -4059
rect -9117 -4161 -9083 -4127
rect -9117 -4229 -9083 -4195
rect -9117 -4297 -9083 -4263
rect -9117 -4365 -9083 -4331
rect -9117 -4433 -9083 -4399
rect -9117 -4513 -9083 -4467
rect -12957 -4547 -12873 -4513
rect -12839 -4547 -12805 -4513
rect -12771 -4547 -12737 -4513
rect -12703 -4547 -12669 -4513
rect -12635 -4547 -12601 -4513
rect -12567 -4547 -12533 -4513
rect -12499 -4547 -12465 -4513
rect -12431 -4547 -12397 -4513
rect -12363 -4547 -12329 -4513
rect -12295 -4547 -12261 -4513
rect -12227 -4547 -12193 -4513
rect -12159 -4547 -12125 -4513
rect -12091 -4547 -12057 -4513
rect -12023 -4547 -11989 -4513
rect -11955 -4547 -11921 -4513
rect -11887 -4547 -11853 -4513
rect -11819 -4547 -11785 -4513
rect -11751 -4547 -11717 -4513
rect -11683 -4547 -11649 -4513
rect -11615 -4547 -11581 -4513
rect -11547 -4547 -11513 -4513
rect -11479 -4547 -11445 -4513
rect -11411 -4547 -11377 -4513
rect -11343 -4547 -11309 -4513
rect -11275 -4547 -11241 -4513
rect -11207 -4547 -11173 -4513
rect -11139 -4547 -11105 -4513
rect -11071 -4547 -11037 -4513
rect -11003 -4547 -10969 -4513
rect -10935 -4547 -10901 -4513
rect -10867 -4547 -10833 -4513
rect -10799 -4547 -10765 -4513
rect -10731 -4547 -10697 -4513
rect -10663 -4547 -10629 -4513
rect -10595 -4547 -10561 -4513
rect -10527 -4547 -10493 -4513
rect -10459 -4547 -10425 -4513
rect -10391 -4547 -10357 -4513
rect -10323 -4547 -10289 -4513
rect -10255 -4547 -10221 -4513
rect -10187 -4547 -10153 -4513
rect -10119 -4547 -10085 -4513
rect -10051 -4547 -10017 -4513
rect -9983 -4547 -9949 -4513
rect -9915 -4547 -9881 -4513
rect -9847 -4547 -9813 -4513
rect -9779 -4547 -9745 -4513
rect -9711 -4547 -9677 -4513
rect -9643 -4547 -9609 -4513
rect -9575 -4547 -9541 -4513
rect -9507 -4547 -9473 -4513
rect -9439 -4547 -9405 -4513
rect -9371 -4547 -9337 -4513
rect -9303 -4547 -9269 -4513
rect -9235 -4547 -9201 -4513
rect -9167 -4547 -9083 -4513
<< viali >>
rect -59 -3057 -45 -3023
rect -45 -3057 -25 -3023
rect 13 -3057 23 -3023
rect 23 -3057 47 -3023
rect 85 -3057 91 -3023
rect 91 -3057 119 -3023
rect 157 -3057 159 -3023
rect 159 -3057 191 -3023
rect 229 -3057 261 -3023
rect 261 -3057 263 -3023
rect 301 -3057 329 -3023
rect 329 -3057 335 -3023
rect 373 -3057 397 -3023
rect 397 -3057 407 -3023
rect 445 -3057 465 -3023
rect 465 -3057 479 -3023
<< metal1 >>
rect 380 140 440 150
rect 140 136 440 140
rect -180 80 -120 90
rect 140 84 384 136
rect 436 84 440 136
rect 140 80 440 84
rect -180 76 100 80
rect -180 24 -176 76
rect -124 24 100 76
rect 380 70 440 80
rect -180 20 100 24
rect -180 10 -120 20
rect 130 -60 280 30
rect -330 -120 280 -60
rect 380 -160 440 -150
rect 140 -164 440 -160
rect -60 -220 0 -210
rect 140 -216 384 -164
rect 436 -216 440 -164
rect 140 -220 440 -216
rect -60 -224 100 -220
rect -60 -276 -56 -224
rect -4 -276 100 -224
rect 380 -230 440 -220
rect -60 -280 100 -276
rect 130 -280 280 -270
rect -60 -290 0 -280
rect 130 -340 520 -280
rect -330 -400 280 -340
rect 380 -460 440 -450
rect 140 -464 440 -460
rect -180 -520 -120 -510
rect 140 -516 384 -464
rect 436 -516 440 -464
rect 140 -520 440 -516
rect -180 -524 100 -520
rect -180 -576 -176 -524
rect -124 -576 100 -524
rect 380 -530 440 -520
rect -180 -580 100 -576
rect 130 -580 180 -570
rect -180 -590 -120 -580
rect 130 -660 280 -580
rect -330 -720 280 -660
rect 380 -760 440 -750
rect 140 -764 440 -760
rect -60 -820 0 -810
rect 140 -816 384 -764
rect 436 -816 440 -764
rect 140 -820 440 -816
rect -60 -824 100 -820
rect -60 -876 -56 -824
rect -4 -876 100 -824
rect 380 -830 440 -820
rect -60 -880 100 -876
rect 130 -880 160 -870
rect -60 -890 0 -880
rect 130 -940 520 -880
rect -330 -1000 280 -940
rect 380 -1060 440 -1050
rect 140 -1064 440 -1060
rect -180 -1120 -120 -1110
rect 140 -1116 384 -1064
rect 436 -1116 440 -1064
rect 140 -1120 440 -1116
rect -180 -1124 100 -1120
rect -180 -1176 -176 -1124
rect -124 -1176 100 -1124
rect 380 -1130 440 -1120
rect -180 -1180 100 -1176
rect -180 -1190 -120 -1180
rect 180 -1260 280 -1180
rect -330 -1320 280 -1260
rect 380 -1360 440 -1350
rect 140 -1364 440 -1360
rect -60 -1420 0 -1410
rect 140 -1416 384 -1364
rect 436 -1416 440 -1364
rect 140 -1420 440 -1416
rect -60 -1424 100 -1420
rect -60 -1476 -56 -1424
rect -4 -1476 100 -1424
rect 380 -1430 440 -1420
rect -60 -1480 100 -1476
rect 130 -1480 200 -1470
rect -60 -1490 0 -1480
rect 130 -1540 520 -1480
rect -330 -1600 280 -1540
rect 380 -1660 440 -1650
rect 140 -1664 440 -1660
rect -60 -1720 0 -1710
rect 140 -1716 384 -1664
rect 436 -1716 440 -1664
rect 140 -1720 440 -1716
rect -60 -1724 100 -1720
rect -60 -1776 -56 -1724
rect -4 -1776 100 -1724
rect 380 -1730 440 -1720
rect -60 -1780 100 -1776
rect 130 -1780 190 -1770
rect -60 -1790 0 -1780
rect 130 -1840 520 -1780
rect -270 -1900 270 -1840
rect 380 -1960 440 -1950
rect 140 -1964 440 -1960
rect -180 -2020 -120 -2010
rect 140 -2016 384 -1964
rect 436 -2016 440 -1964
rect 140 -2020 440 -2016
rect -180 -2024 100 -2020
rect -180 -2076 -176 -2024
rect -124 -2076 100 -2024
rect 380 -2030 440 -2020
rect -180 -2080 100 -2076
rect -180 -2090 -120 -2080
rect 140 -2160 260 -2080
rect -330 -2220 260 -2160
rect 380 -2260 440 -2250
rect 140 -2264 440 -2260
rect -180 -2320 -120 -2310
rect 140 -2316 384 -2264
rect 436 -2316 440 -2264
rect 140 -2320 440 -2316
rect -180 -2324 100 -2320
rect -180 -2376 -176 -2324
rect -124 -2376 100 -2324
rect 380 -2330 440 -2320
rect -180 -2380 100 -2376
rect -180 -2390 -120 -2380
rect 140 -2460 280 -2380
rect -330 -2520 280 -2460
rect 380 -2560 440 -2550
rect 140 -2564 440 -2560
rect -60 -2620 0 -2610
rect 140 -2616 384 -2564
rect 436 -2616 440 -2564
rect 140 -2620 440 -2616
rect -60 -2624 100 -2620
rect -60 -2676 -56 -2624
rect -4 -2676 100 -2624
rect 380 -2630 440 -2620
rect -60 -2680 100 -2676
rect -60 -2690 0 -2680
rect 200 -2960 260 -2680
rect -100 -3023 560 -3000
rect -100 -3057 -59 -3023
rect -25 -3057 13 -3023
rect 47 -3057 85 -3023
rect 119 -3057 157 -3023
rect 191 -3057 229 -3023
rect 263 -3057 301 -3023
rect 335 -3057 373 -3023
rect 407 -3057 445 -3023
rect 479 -3057 560 -3023
rect -100 -3080 560 -3057
<< via1 >>
rect 384 84 436 136
rect -176 24 -124 76
rect 384 -216 436 -164
rect -56 -276 -4 -224
rect 384 -516 436 -464
rect -176 -576 -124 -524
rect 384 -816 436 -764
rect -56 -876 -4 -824
rect 384 -1116 436 -1064
rect -176 -1176 -124 -1124
rect 384 -1416 436 -1364
rect -56 -1476 -4 -1424
rect 384 -1716 436 -1664
rect -56 -1776 -4 -1724
rect 384 -2016 436 -1964
rect -176 -2076 -124 -2024
rect 384 -2316 436 -2264
rect -176 -2376 -124 -2324
rect 384 -2616 436 -2564
rect -56 -2676 -4 -2624
<< metal2 >>
rect -180 80 -120 240
rect -180 76 -110 80
rect -180 24 -176 76
rect -124 24 -110 76
rect -180 20 -110 24
rect -180 -520 -120 20
rect -60 -220 0 240
rect 370 136 450 140
rect 370 84 384 136
rect 436 84 450 136
rect 370 80 450 84
rect 380 -150 440 80
rect 380 -160 460 -150
rect 370 -162 460 -160
rect 370 -164 392 -162
rect 370 -216 384 -164
rect 370 -218 392 -216
rect 448 -218 460 -162
rect 370 -220 460 -218
rect -70 -224 10 -220
rect -70 -276 -56 -224
rect -4 -276 10 -224
rect 380 -230 460 -220
rect -70 -280 10 -276
rect -180 -524 -110 -520
rect -180 -576 -176 -524
rect -124 -576 -110 -524
rect -180 -580 -110 -576
rect -180 -1120 -120 -580
rect -60 -820 0 -280
rect 370 -464 450 -460
rect 370 -516 384 -464
rect 436 -516 450 -464
rect 370 -520 450 -516
rect 380 -750 440 -520
rect 380 -760 460 -750
rect 370 -762 460 -760
rect 370 -764 392 -762
rect 370 -816 384 -764
rect 370 -818 392 -816
rect 448 -818 460 -762
rect 370 -820 460 -818
rect -70 -824 10 -820
rect -70 -876 -56 -824
rect -4 -876 10 -824
rect 380 -830 460 -820
rect -70 -880 10 -876
rect -180 -1124 -110 -1120
rect -180 -1176 -176 -1124
rect -124 -1176 -110 -1124
rect -180 -1180 -110 -1176
rect -180 -2020 -120 -1180
rect -60 -1420 0 -880
rect 370 -1064 450 -1060
rect 370 -1116 384 -1064
rect 436 -1116 450 -1064
rect 370 -1120 450 -1116
rect 380 -1350 440 -1120
rect 380 -1360 460 -1350
rect 370 -1362 460 -1360
rect 370 -1364 392 -1362
rect 370 -1416 384 -1364
rect 370 -1418 392 -1416
rect 448 -1418 460 -1362
rect 370 -1420 460 -1418
rect -70 -1424 10 -1420
rect -70 -1476 -56 -1424
rect -4 -1476 10 -1424
rect 380 -1430 460 -1420
rect -70 -1480 10 -1476
rect -60 -1720 0 -1480
rect 370 -1664 450 -1660
rect 370 -1716 384 -1664
rect 436 -1716 450 -1664
rect 370 -1720 450 -1716
rect -70 -1724 10 -1720
rect -70 -1776 -56 -1724
rect -4 -1776 10 -1724
rect -70 -1780 10 -1776
rect -180 -2024 -110 -2020
rect -180 -2076 -176 -2024
rect -124 -2076 -110 -2024
rect -180 -2080 -110 -2076
rect -180 -2320 -120 -2080
rect -180 -2324 -110 -2320
rect -180 -2376 -176 -2324
rect -124 -2376 -110 -2324
rect -180 -2380 -110 -2376
rect -180 -2980 -120 -2380
rect -60 -2620 0 -1780
rect 380 -1950 440 -1720
rect 380 -1960 460 -1950
rect 370 -1962 460 -1960
rect 370 -1964 392 -1962
rect 370 -2016 384 -1964
rect 370 -2018 392 -2016
rect 448 -2018 460 -1962
rect 370 -2020 460 -2018
rect 380 -2030 460 -2020
rect 370 -2264 450 -2260
rect 370 -2316 384 -2264
rect 436 -2316 450 -2264
rect 370 -2320 450 -2316
rect 380 -2550 440 -2320
rect 380 -2560 460 -2550
rect 370 -2562 460 -2560
rect 370 -2564 392 -2562
rect 370 -2616 384 -2564
rect 370 -2618 392 -2616
rect 448 -2618 460 -2562
rect 370 -2620 460 -2618
rect -70 -2624 10 -2620
rect -70 -2676 -56 -2624
rect -4 -2676 10 -2624
rect 380 -2630 460 -2620
rect -70 -2680 10 -2676
rect -60 -2980 0 -2680
<< via2 >>
rect 392 -164 448 -162
rect 392 -216 436 -164
rect 436 -216 448 -164
rect 392 -218 448 -216
rect 392 -764 448 -762
rect 392 -816 436 -764
rect 436 -816 448 -764
rect 392 -818 448 -816
rect 392 -1364 448 -1362
rect 392 -1416 436 -1364
rect 436 -1416 448 -1364
rect 392 -1418 448 -1416
rect 392 -1964 448 -1962
rect 392 -2016 436 -1964
rect 436 -2016 448 -1964
rect 392 -2018 448 -2016
rect 392 -2564 448 -2562
rect 392 -2616 436 -2564
rect 436 -2616 448 -2564
rect 392 -2618 448 -2616
<< metal3 >>
rect 870 -108 990 -90
rect 870 -150 898 -108
rect 380 -162 898 -150
rect 380 -218 392 -162
rect 448 -172 898 -162
rect 962 -172 990 -108
rect 448 -218 990 -172
rect 380 -228 990 -218
rect 380 -230 898 -228
rect 870 -292 898 -230
rect 962 -292 990 -228
rect 870 -310 990 -292
rect 1050 -718 1170 -700
rect 1050 -750 1078 -718
rect 380 -762 1078 -750
rect 380 -818 392 -762
rect 448 -782 1078 -762
rect 1142 -782 1170 -718
rect 448 -818 1170 -782
rect 380 -830 1170 -818
rect 1050 -838 1170 -830
rect 1050 -902 1078 -838
rect 1142 -902 1170 -838
rect 1050 -920 1170 -902
rect 1240 -1308 1360 -1290
rect 1240 -1350 1268 -1308
rect 380 -1362 1268 -1350
rect 380 -1418 392 -1362
rect 448 -1372 1268 -1362
rect 1332 -1372 1360 -1308
rect 448 -1418 1360 -1372
rect 380 -1428 1360 -1418
rect 380 -1430 1268 -1428
rect 1240 -1492 1268 -1430
rect 1332 -1492 1360 -1428
rect 1240 -1510 1360 -1492
rect 1420 -1888 1540 -1870
rect 1420 -1950 1448 -1888
rect 380 -1952 1448 -1950
rect 1512 -1952 1540 -1888
rect 380 -1962 1540 -1952
rect 380 -2018 392 -1962
rect 448 -2008 1540 -1962
rect 448 -2018 1448 -2008
rect 380 -2030 1448 -2018
rect 1420 -2072 1448 -2030
rect 1512 -2072 1540 -2008
rect 1420 -2090 1540 -2072
rect 380 -2562 690 -2550
rect 380 -2618 392 -2562
rect 448 -2618 690 -2562
rect 380 -2630 690 -2618
<< via3 >>
rect 898 -172 962 -108
rect 898 -292 962 -228
rect 1078 -782 1142 -718
rect 1078 -902 1142 -838
rect 1268 -1372 1332 -1308
rect 1268 -1492 1332 -1428
rect 1448 -1952 1512 -1888
rect 1448 -2072 1512 -2008
<< metal4 >>
rect 870 -108 990 -90
rect 870 -172 898 -108
rect 962 -172 990 -108
rect 870 -228 990 -172
rect 870 -292 898 -228
rect 962 -292 990 -228
rect 870 -310 990 -292
rect 1050 -718 1170 -700
rect 1050 -782 1078 -718
rect 1142 -782 1170 -718
rect 1050 -838 1170 -782
rect 1050 -902 1078 -838
rect 1142 -902 1170 -838
rect 1050 -920 1170 -902
rect 1240 -1308 1360 -1290
rect 1240 -1372 1268 -1308
rect 1332 -1372 1360 -1308
rect 1240 -1428 1360 -1372
rect 1240 -1492 1268 -1428
rect 1332 -1492 1360 -1428
rect 1240 -1510 1360 -1492
rect 1420 -1888 1540 -1870
rect 1420 -1952 1448 -1888
rect 1512 -1952 1540 -1888
rect 1420 -2008 1540 -1952
rect 1420 -2072 1448 -2008
rect 1512 -2072 1540 -2008
rect 1420 -2090 1540 -2072
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_0
timestamp 1757161594
transform 0 -1 203 1 0 -2347
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_1
timestamp 1757161594
transform 0 -1 203 1 0 -2647
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_2
timestamp 1757161594
transform 0 -1 203 1 0 -1747
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_3
timestamp 1757161594
transform 0 -1 203 1 0 -2047
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_4
timestamp 1757161594
transform 0 -1 203 1 0 -1447
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_5
timestamp 1757161594
transform 0 -1 203 1 0 -847
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_6
timestamp 1757161594
transform 0 -1 203 1 0 -1147
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_7
timestamp 1757161594
transform 0 -1 203 1 0 -247
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_8
timestamp 1757161594
transform 0 -1 203 1 0 -547
box -99 -157 99 157
use sky130_fd_pr__nfet_01v8_lvt_6DE3T6  sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9
timestamp 1757161594
transform 0 -1 203 1 0 53
box -99 -157 99 157
<< labels >>
rlabel metal2 s -60 -2980 0 -2920 4 en_1
port 1 nsew
rlabel metal2 s -180 -2980 -120 -2920 4 en_2
port 2 nsew
rlabel metal1 s 200 -2960 260 -2900 4 beta
port 3 nsew
rlabel metal1 s 460 -1840 520 -1780 4 Vbias1
port 4 nsew
rlabel metal1 s 460 -1540 520 -1480 4 Vbias2
port 5 nsew
rlabel metal1 s 460 -940 520 -880 4 Vbias3
port 6 nsew
rlabel metal1 s 460 -340 520 -280 4 Vbias4
port 7 nsew
<< end >>
