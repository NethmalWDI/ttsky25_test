magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -2084 -107 2084 45
<< nmoslvt >>
rect -2000 -81 2000 19
<< ndiff >>
rect -2058 -14 -2000 19
rect -2058 -48 -2046 -14
rect -2012 -48 -2000 -14
rect -2058 -81 -2000 -48
rect 2000 -14 2058 19
rect 2000 -48 2012 -14
rect 2046 -48 2058 -14
rect 2000 -81 2058 -48
<< ndiffc >>
rect -2046 -48 -2012 -14
rect 2012 -48 2046 -14
<< poly >>
rect -2000 91 2000 107
rect -2000 57 -1955 91
rect -1921 57 -1887 91
rect -1853 57 -1819 91
rect -1785 57 -1751 91
rect -1717 57 -1683 91
rect -1649 57 -1615 91
rect -1581 57 -1547 91
rect -1513 57 -1479 91
rect -1445 57 -1411 91
rect -1377 57 -1343 91
rect -1309 57 -1275 91
rect -1241 57 -1207 91
rect -1173 57 -1139 91
rect -1105 57 -1071 91
rect -1037 57 -1003 91
rect -969 57 -935 91
rect -901 57 -867 91
rect -833 57 -799 91
rect -765 57 -731 91
rect -697 57 -663 91
rect -629 57 -595 91
rect -561 57 -527 91
rect -493 57 -459 91
rect -425 57 -391 91
rect -357 57 -323 91
rect -289 57 -255 91
rect -221 57 -187 91
rect -153 57 -119 91
rect -85 57 -51 91
rect -17 57 17 91
rect 51 57 85 91
rect 119 57 153 91
rect 187 57 221 91
rect 255 57 289 91
rect 323 57 357 91
rect 391 57 425 91
rect 459 57 493 91
rect 527 57 561 91
rect 595 57 629 91
rect 663 57 697 91
rect 731 57 765 91
rect 799 57 833 91
rect 867 57 901 91
rect 935 57 969 91
rect 1003 57 1037 91
rect 1071 57 1105 91
rect 1139 57 1173 91
rect 1207 57 1241 91
rect 1275 57 1309 91
rect 1343 57 1377 91
rect 1411 57 1445 91
rect 1479 57 1513 91
rect 1547 57 1581 91
rect 1615 57 1649 91
rect 1683 57 1717 91
rect 1751 57 1785 91
rect 1819 57 1853 91
rect 1887 57 1921 91
rect 1955 57 2000 91
rect -2000 19 2000 57
rect -2000 -107 2000 -81
<< polycont >>
rect -1955 57 -1921 91
rect -1887 57 -1853 91
rect -1819 57 -1785 91
rect -1751 57 -1717 91
rect -1683 57 -1649 91
rect -1615 57 -1581 91
rect -1547 57 -1513 91
rect -1479 57 -1445 91
rect -1411 57 -1377 91
rect -1343 57 -1309 91
rect -1275 57 -1241 91
rect -1207 57 -1173 91
rect -1139 57 -1105 91
rect -1071 57 -1037 91
rect -1003 57 -969 91
rect -935 57 -901 91
rect -867 57 -833 91
rect -799 57 -765 91
rect -731 57 -697 91
rect -663 57 -629 91
rect -595 57 -561 91
rect -527 57 -493 91
rect -459 57 -425 91
rect -391 57 -357 91
rect -323 57 -289 91
rect -255 57 -221 91
rect -187 57 -153 91
rect -119 57 -85 91
rect -51 57 -17 91
rect 17 57 51 91
rect 85 57 119 91
rect 153 57 187 91
rect 221 57 255 91
rect 289 57 323 91
rect 357 57 391 91
rect 425 57 459 91
rect 493 57 527 91
rect 561 57 595 91
rect 629 57 663 91
rect 697 57 731 91
rect 765 57 799 91
rect 833 57 867 91
rect 901 57 935 91
rect 969 57 1003 91
rect 1037 57 1071 91
rect 1105 57 1139 91
rect 1173 57 1207 91
rect 1241 57 1275 91
rect 1309 57 1343 91
rect 1377 57 1411 91
rect 1445 57 1479 91
rect 1513 57 1547 91
rect 1581 57 1615 91
rect 1649 57 1683 91
rect 1717 57 1751 91
rect 1785 57 1819 91
rect 1853 57 1887 91
rect 1921 57 1955 91
<< locali >>
rect -2000 57 -1961 91
rect -1921 57 -1889 91
rect -1853 57 -1819 91
rect -1783 57 -1751 91
rect -1711 57 -1683 91
rect -1639 57 -1615 91
rect -1567 57 -1547 91
rect -1495 57 -1479 91
rect -1423 57 -1411 91
rect -1351 57 -1343 91
rect -1279 57 -1275 91
rect -1173 57 -1169 91
rect -1105 57 -1097 91
rect -1037 57 -1025 91
rect -969 57 -953 91
rect -901 57 -881 91
rect -833 57 -809 91
rect -765 57 -737 91
rect -697 57 -665 91
rect -629 57 -595 91
rect -559 57 -527 91
rect -487 57 -459 91
rect -415 57 -391 91
rect -343 57 -323 91
rect -271 57 -255 91
rect -199 57 -187 91
rect -127 57 -119 91
rect -55 57 -51 91
rect 51 57 55 91
rect 119 57 127 91
rect 187 57 199 91
rect 255 57 271 91
rect 323 57 343 91
rect 391 57 415 91
rect 459 57 487 91
rect 527 57 559 91
rect 595 57 629 91
rect 665 57 697 91
rect 737 57 765 91
rect 809 57 833 91
rect 881 57 901 91
rect 953 57 969 91
rect 1025 57 1037 91
rect 1097 57 1105 91
rect 1169 57 1173 91
rect 1275 57 1279 91
rect 1343 57 1351 91
rect 1411 57 1423 91
rect 1479 57 1495 91
rect 1547 57 1567 91
rect 1615 57 1639 91
rect 1683 57 1711 91
rect 1751 57 1783 91
rect 1819 57 1853 91
rect 1889 57 1921 91
rect 1961 57 2000 91
rect -2046 -14 -2012 23
rect -2046 -85 -2012 -48
rect 2012 -14 2046 23
rect 2012 -85 2046 -48
<< viali >>
rect -1961 57 -1955 91
rect -1955 57 -1927 91
rect -1889 57 -1887 91
rect -1887 57 -1855 91
rect -1817 57 -1785 91
rect -1785 57 -1783 91
rect -1745 57 -1717 91
rect -1717 57 -1711 91
rect -1673 57 -1649 91
rect -1649 57 -1639 91
rect -1601 57 -1581 91
rect -1581 57 -1567 91
rect -1529 57 -1513 91
rect -1513 57 -1495 91
rect -1457 57 -1445 91
rect -1445 57 -1423 91
rect -1385 57 -1377 91
rect -1377 57 -1351 91
rect -1313 57 -1309 91
rect -1309 57 -1279 91
rect -1241 57 -1207 91
rect -1169 57 -1139 91
rect -1139 57 -1135 91
rect -1097 57 -1071 91
rect -1071 57 -1063 91
rect -1025 57 -1003 91
rect -1003 57 -991 91
rect -953 57 -935 91
rect -935 57 -919 91
rect -881 57 -867 91
rect -867 57 -847 91
rect -809 57 -799 91
rect -799 57 -775 91
rect -737 57 -731 91
rect -731 57 -703 91
rect -665 57 -663 91
rect -663 57 -631 91
rect -593 57 -561 91
rect -561 57 -559 91
rect -521 57 -493 91
rect -493 57 -487 91
rect -449 57 -425 91
rect -425 57 -415 91
rect -377 57 -357 91
rect -357 57 -343 91
rect -305 57 -289 91
rect -289 57 -271 91
rect -233 57 -221 91
rect -221 57 -199 91
rect -161 57 -153 91
rect -153 57 -127 91
rect -89 57 -85 91
rect -85 57 -55 91
rect -17 57 17 91
rect 55 57 85 91
rect 85 57 89 91
rect 127 57 153 91
rect 153 57 161 91
rect 199 57 221 91
rect 221 57 233 91
rect 271 57 289 91
rect 289 57 305 91
rect 343 57 357 91
rect 357 57 377 91
rect 415 57 425 91
rect 425 57 449 91
rect 487 57 493 91
rect 493 57 521 91
rect 559 57 561 91
rect 561 57 593 91
rect 631 57 663 91
rect 663 57 665 91
rect 703 57 731 91
rect 731 57 737 91
rect 775 57 799 91
rect 799 57 809 91
rect 847 57 867 91
rect 867 57 881 91
rect 919 57 935 91
rect 935 57 953 91
rect 991 57 1003 91
rect 1003 57 1025 91
rect 1063 57 1071 91
rect 1071 57 1097 91
rect 1135 57 1139 91
rect 1139 57 1169 91
rect 1207 57 1241 91
rect 1279 57 1309 91
rect 1309 57 1313 91
rect 1351 57 1377 91
rect 1377 57 1385 91
rect 1423 57 1445 91
rect 1445 57 1457 91
rect 1495 57 1513 91
rect 1513 57 1529 91
rect 1567 57 1581 91
rect 1581 57 1601 91
rect 1639 57 1649 91
rect 1649 57 1673 91
rect 1711 57 1717 91
rect 1717 57 1745 91
rect 1783 57 1785 91
rect 1785 57 1817 91
rect 1855 57 1887 91
rect 1887 57 1889 91
rect 1927 57 1955 91
rect 1955 57 1961 91
rect -2046 -48 -2012 -14
rect 2012 -48 2046 -14
<< metal1 >>
rect -1996 91 1996 97
rect -1996 57 -1961 91
rect -1927 57 -1889 91
rect -1855 57 -1817 91
rect -1783 57 -1745 91
rect -1711 57 -1673 91
rect -1639 57 -1601 91
rect -1567 57 -1529 91
rect -1495 57 -1457 91
rect -1423 57 -1385 91
rect -1351 57 -1313 91
rect -1279 57 -1241 91
rect -1207 57 -1169 91
rect -1135 57 -1097 91
rect -1063 57 -1025 91
rect -991 57 -953 91
rect -919 57 -881 91
rect -847 57 -809 91
rect -775 57 -737 91
rect -703 57 -665 91
rect -631 57 -593 91
rect -559 57 -521 91
rect -487 57 -449 91
rect -415 57 -377 91
rect -343 57 -305 91
rect -271 57 -233 91
rect -199 57 -161 91
rect -127 57 -89 91
rect -55 57 -17 91
rect 17 57 55 91
rect 89 57 127 91
rect 161 57 199 91
rect 233 57 271 91
rect 305 57 343 91
rect 377 57 415 91
rect 449 57 487 91
rect 521 57 559 91
rect 593 57 631 91
rect 665 57 703 91
rect 737 57 775 91
rect 809 57 847 91
rect 881 57 919 91
rect 953 57 991 91
rect 1025 57 1063 91
rect 1097 57 1135 91
rect 1169 57 1207 91
rect 1241 57 1279 91
rect 1313 57 1351 91
rect 1385 57 1423 91
rect 1457 57 1495 91
rect 1529 57 1567 91
rect 1601 57 1639 91
rect 1673 57 1711 91
rect 1745 57 1783 91
rect 1817 57 1855 91
rect 1889 57 1927 91
rect 1961 57 1996 91
rect -1996 51 1996 57
rect -2052 -14 -2006 19
rect -2052 -48 -2046 -14
rect -2012 -48 -2006 -14
rect -2052 -81 -2006 -48
rect 2006 -14 2052 19
rect 2006 -48 2012 -14
rect 2046 -48 2052 -14
rect 2006 -81 2052 -48
<< end >>
