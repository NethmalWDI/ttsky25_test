magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -500 -2860 2080 2840
<< nsubdiff >>
rect -460 2777 1980 2800
rect -460 2743 -359 2777
rect -325 2743 -291 2777
rect -257 2743 -223 2777
rect -189 2743 -155 2777
rect -121 2743 -87 2777
rect -53 2743 -19 2777
rect 15 2743 49 2777
rect 83 2743 117 2777
rect 151 2743 185 2777
rect 219 2743 253 2777
rect 287 2743 321 2777
rect 355 2743 389 2777
rect 423 2743 457 2777
rect 491 2743 525 2777
rect 559 2743 593 2777
rect 627 2743 661 2777
rect 695 2743 729 2777
rect 763 2743 797 2777
rect 831 2743 865 2777
rect 899 2743 933 2777
rect 967 2743 1001 2777
rect 1035 2743 1069 2777
rect 1103 2743 1137 2777
rect 1171 2743 1205 2777
rect 1239 2743 1273 2777
rect 1307 2743 1341 2777
rect 1375 2743 1409 2777
rect 1443 2743 1477 2777
rect 1511 2743 1545 2777
rect 1579 2743 1613 2777
rect 1647 2743 1681 2777
rect 1715 2743 1749 2777
rect 1783 2743 1817 2777
rect 1851 2743 1885 2777
rect 1919 2743 1980 2777
rect -460 2720 1980 2743
rect -460 -2780 -420 2720
rect 1940 -2780 1980 2720
rect -460 -2820 1980 -2780
<< nsubdiffcont >>
rect -359 2743 -325 2777
rect -291 2743 -257 2777
rect -223 2743 -189 2777
rect -155 2743 -121 2777
rect -87 2743 -53 2777
rect -19 2743 15 2777
rect 49 2743 83 2777
rect 117 2743 151 2777
rect 185 2743 219 2777
rect 253 2743 287 2777
rect 321 2743 355 2777
rect 389 2743 423 2777
rect 457 2743 491 2777
rect 525 2743 559 2777
rect 593 2743 627 2777
rect 661 2743 695 2777
rect 729 2743 763 2777
rect 797 2743 831 2777
rect 865 2743 899 2777
rect 933 2743 967 2777
rect 1001 2743 1035 2777
rect 1069 2743 1103 2777
rect 1137 2743 1171 2777
rect 1205 2743 1239 2777
rect 1273 2743 1307 2777
rect 1341 2743 1375 2777
rect 1409 2743 1443 2777
rect 1477 2743 1511 2777
rect 1545 2743 1579 2777
rect 1613 2743 1647 2777
rect 1681 2743 1715 2777
rect 1749 2743 1783 2777
rect 1817 2743 1851 2777
rect 1885 2743 1919 2777
<< locali >>
rect -460 2777 1980 2800
rect -460 2743 -359 2777
rect -319 2743 -291 2777
rect -247 2743 -223 2777
rect -175 2743 -155 2777
rect -103 2743 -87 2777
rect -31 2743 -19 2777
rect 41 2743 49 2777
rect 113 2743 117 2777
rect 219 2743 223 2777
rect 287 2743 295 2777
rect 355 2743 367 2777
rect 423 2743 439 2777
rect 491 2743 511 2777
rect 559 2743 583 2777
rect 627 2743 655 2777
rect 695 2743 727 2777
rect 763 2743 797 2777
rect 833 2743 865 2777
rect 905 2743 933 2777
rect 977 2743 1001 2777
rect 1049 2743 1069 2777
rect 1121 2743 1137 2777
rect 1193 2743 1205 2777
rect 1265 2743 1273 2777
rect 1337 2743 1341 2777
rect 1443 2743 1447 2777
rect 1511 2743 1519 2777
rect 1579 2743 1591 2777
rect 1647 2743 1663 2777
rect 1715 2743 1735 2777
rect 1783 2743 1807 2777
rect 1851 2743 1879 2777
rect 1919 2743 1980 2777
rect -460 2720 1980 2743
rect -460 -2780 -420 2720
rect 1940 -2780 1980 2720
rect -460 -2820 1980 -2780
<< viali >>
rect -353 2743 -325 2777
rect -325 2743 -319 2777
rect -281 2743 -257 2777
rect -257 2743 -247 2777
rect -209 2743 -189 2777
rect -189 2743 -175 2777
rect -137 2743 -121 2777
rect -121 2743 -103 2777
rect -65 2743 -53 2777
rect -53 2743 -31 2777
rect 7 2743 15 2777
rect 15 2743 41 2777
rect 79 2743 83 2777
rect 83 2743 113 2777
rect 151 2743 185 2777
rect 223 2743 253 2777
rect 253 2743 257 2777
rect 295 2743 321 2777
rect 321 2743 329 2777
rect 367 2743 389 2777
rect 389 2743 401 2777
rect 439 2743 457 2777
rect 457 2743 473 2777
rect 511 2743 525 2777
rect 525 2743 545 2777
rect 583 2743 593 2777
rect 593 2743 617 2777
rect 655 2743 661 2777
rect 661 2743 689 2777
rect 727 2743 729 2777
rect 729 2743 761 2777
rect 799 2743 831 2777
rect 831 2743 833 2777
rect 871 2743 899 2777
rect 899 2743 905 2777
rect 943 2743 967 2777
rect 967 2743 977 2777
rect 1015 2743 1035 2777
rect 1035 2743 1049 2777
rect 1087 2743 1103 2777
rect 1103 2743 1121 2777
rect 1159 2743 1171 2777
rect 1171 2743 1193 2777
rect 1231 2743 1239 2777
rect 1239 2743 1265 2777
rect 1303 2743 1307 2777
rect 1307 2743 1337 2777
rect 1375 2743 1409 2777
rect 1447 2743 1477 2777
rect 1477 2743 1481 2777
rect 1519 2743 1545 2777
rect 1545 2743 1553 2777
rect 1591 2743 1613 2777
rect 1613 2743 1625 2777
rect 1663 2743 1681 2777
rect 1681 2743 1697 2777
rect 1735 2743 1749 2777
rect 1749 2743 1769 2777
rect 1807 2743 1817 2777
rect 1817 2743 1841 2777
rect 1879 2743 1885 2777
rect 1885 2743 1913 2777
<< metal1 >>
rect -460 2777 1980 2800
rect -460 2743 -353 2777
rect -319 2743 -281 2777
rect -247 2743 -209 2777
rect -175 2743 -137 2777
rect -103 2743 -65 2777
rect -31 2743 7 2777
rect 41 2743 79 2777
rect 113 2743 151 2777
rect 185 2743 223 2777
rect 257 2743 295 2777
rect 329 2743 367 2777
rect 401 2743 439 2777
rect 473 2743 511 2777
rect 545 2743 583 2777
rect 617 2743 655 2777
rect 689 2743 727 2777
rect 761 2743 799 2777
rect 833 2743 871 2777
rect 905 2743 943 2777
rect 977 2743 1015 2777
rect 1049 2743 1087 2777
rect 1121 2743 1159 2777
rect 1193 2743 1231 2777
rect 1265 2743 1303 2777
rect 1337 2743 1375 2777
rect 1409 2743 1447 2777
rect 1481 2743 1519 2777
rect 1553 2743 1591 2777
rect 1625 2743 1663 2777
rect 1697 2743 1735 2777
rect 1769 2743 1807 2777
rect 1841 2743 1879 2777
rect 1913 2743 1980 2777
rect -460 2720 1980 2743
rect -200 2660 -120 2720
rect -340 2600 1900 2660
rect -200 2500 -120 2600
rect 200 2500 260 2600
rect 600 2500 660 2600
rect 1000 2500 1060 2600
rect 1400 2500 1480 2600
rect 1800 2500 1900 2600
rect -340 2440 -120 2500
rect 60 2440 260 2500
rect 460 2440 660 2500
rect 860 2440 1060 2500
rect 1260 2440 1480 2500
rect 1660 2440 1900 2500
rect -200 2360 -120 2440
rect -340 2300 -120 2360
rect 472 2365 558 2366
rect 64 2357 150 2358
rect 64 2305 81 2357
rect 133 2305 150 2357
rect 472 2313 489 2365
rect 541 2313 558 2365
rect 1268 2363 1354 2364
rect 873 2355 959 2356
rect 873 2303 890 2355
rect 942 2303 959 2355
rect 1268 2311 1285 2363
rect 1337 2311 1354 2363
rect 1800 2360 1900 2440
rect 1660 2300 1900 2360
rect -200 300 -120 2300
rect -570 220 -490 300
rect -450 296 -370 300
rect -450 244 -436 296
rect -384 244 -370 296
rect -450 -2284 -370 244
rect -340 240 -120 300
rect -200 -200 -120 240
rect 62 291 148 292
rect 62 239 79 291
rect 131 239 148 291
rect 200 -63 280 2240
rect 460 177 540 300
rect 456 176 542 177
rect 456 124 473 176
rect 525 124 542 176
rect 460 120 540 124
rect 600 57 680 2240
rect 860 179 940 300
rect 856 178 942 179
rect 856 126 873 178
rect 925 126 942 178
rect 860 120 940 126
rect 1000 58 1080 2240
rect 1264 288 1350 289
rect 1264 236 1281 288
rect 1333 236 1350 288
rect 995 57 1081 58
rect 598 56 684 57
rect 598 4 615 56
rect 667 4 684 56
rect 995 5 1012 57
rect 1064 5 1081 57
rect 193 -64 280 -63
rect 193 -116 210 -64
rect 262 -116 280 -64
rect -340 -260 -120 -200
rect 51 -201 137 -200
rect 51 -253 68 -201
rect 120 -253 137 -201
rect -200 -2260 -120 -260
rect 200 -2220 280 -116
rect 461 -201 547 -200
rect 461 -253 478 -201
rect 530 -253 547 -201
rect 600 -2220 680 4
rect 858 -203 944 -202
rect 858 -255 875 -203
rect 927 -255 944 -203
rect 1000 -2220 1080 5
rect 1400 -64 1480 2240
rect 1800 2200 1900 2300
rect 1820 300 1900 2200
rect 1660 240 1900 300
rect 1397 -65 1483 -64
rect 1397 -117 1414 -65
rect 1466 -117 1483 -65
rect 1260 -201 1346 -200
rect 1260 -253 1277 -201
rect 1329 -253 1346 -201
rect 1400 -2220 1480 -117
rect 1820 -180 1900 240
rect 1660 -260 1900 -180
rect 1800 -320 1900 -260
rect 1820 -2180 1900 -320
rect 1800 -2260 1900 -2180
rect -450 -2336 -436 -2284
rect -384 -2336 -370 -2284
rect -320 -2320 -120 -2260
rect 1261 -2276 1347 -2275
rect -450 -2340 -370 -2336
rect -200 -2500 -120 -2320
rect 62 -2278 148 -2277
rect 62 -2330 79 -2278
rect 131 -2330 148 -2278
rect 460 -2403 560 -2280
rect 460 -2455 482 -2403
rect 534 -2455 560 -2403
rect 460 -2460 560 -2455
rect 860 -2400 960 -2280
rect 1261 -2328 1278 -2276
rect 1330 -2328 1347 -2276
rect 1660 -2320 1900 -2260
rect 860 -2452 881 -2400
rect 933 -2452 960 -2400
rect 860 -2460 960 -2452
rect 1800 -2500 1900 -2320
rect 2000 176 2080 180
rect 2000 124 2014 176
rect 2066 124 2080 176
rect 2000 -2402 2080 124
rect 1996 -2403 2080 -2402
rect 1996 -2455 2013 -2403
rect 2065 -2455 2080 -2403
rect 2000 -2460 2080 -2455
rect -340 -2560 -120 -2500
rect 60 -2560 260 -2520
rect 460 -2560 660 -2520
rect 860 -2560 1060 -2520
rect 1260 -2560 1460 -2500
rect 1660 -2560 1900 -2500
rect -200 -2660 -120 -2560
rect 200 -2660 260 -2560
rect 580 -2660 660 -2560
rect 1000 -2660 1060 -2560
rect 1400 -2660 1460 -2560
rect 1800 -2660 1900 -2560
rect -340 -2720 1900 -2660
<< via1 >>
rect 81 2305 133 2357
rect 489 2313 541 2365
rect 890 2303 942 2355
rect 1285 2311 1337 2363
rect -436 244 -384 296
rect 79 239 131 291
rect 473 124 525 176
rect 873 126 925 178
rect 1281 236 1333 288
rect 615 4 667 56
rect 1012 5 1064 57
rect 210 -116 262 -64
rect 68 -253 120 -201
rect 478 -253 530 -201
rect 875 -255 927 -203
rect 1414 -117 1466 -65
rect 1277 -253 1329 -201
rect -436 -2336 -384 -2284
rect 79 -2330 131 -2278
rect 482 -2455 534 -2403
rect 1278 -2328 1330 -2276
rect 881 -2452 933 -2400
rect 2014 124 2066 176
rect 2013 -2455 2065 -2403
<< metal2 >>
rect -340 2368 1980 2380
rect -340 2365 1912 2368
rect -340 2357 489 2365
rect -340 2305 81 2357
rect 133 2313 489 2357
rect 541 2363 1912 2365
rect 541 2355 1285 2363
rect 541 2313 890 2355
rect 133 2305 890 2313
rect -340 2303 890 2305
rect 942 2311 1285 2355
rect 1337 2312 1912 2363
rect 1968 2312 1980 2368
rect 1337 2311 1980 2312
rect 942 2303 1980 2311
rect -340 2300 1980 2303
rect 74 2295 140 2300
rect 883 2293 949 2300
rect 72 300 138 302
rect -570 296 1360 300
rect -570 244 -436 296
rect -384 291 1360 296
rect -384 244 79 291
rect -570 240 79 244
rect -570 220 -490 240
rect 72 239 79 240
rect 131 288 1360 291
rect 131 240 1281 288
rect 131 239 138 240
rect 72 229 138 239
rect 1274 236 1281 240
rect 1333 240 1360 288
rect 1333 236 1340 240
rect 1274 226 1340 236
rect 466 180 532 187
rect 866 180 932 189
rect -570 178 2080 180
rect -570 176 873 178
rect -570 124 473 176
rect 525 126 873 176
rect 925 176 2080 178
rect 925 126 2014 176
rect 525 124 2014 126
rect 2066 124 2080 176
rect -570 120 2080 124
rect 466 114 532 120
rect 866 116 932 120
rect 1050 68 1250 70
rect 608 60 674 67
rect 1005 60 1250 68
rect 600 58 1250 60
rect 600 57 1092 58
rect 600 56 1012 57
rect 600 4 615 56
rect 667 5 1012 56
rect 1064 5 1092 57
rect 667 4 1092 5
rect 600 2 1092 4
rect 1148 2 1182 58
rect 1238 2 1250 58
rect 600 0 1250 2
rect 608 -6 674 0
rect 1005 -5 1250 0
rect 1050 -10 1250 -5
rect 203 -60 269 -53
rect 1407 -60 1473 -54
rect -450 -64 1480 -60
rect -450 -72 210 -64
rect -450 -128 -438 -72
rect -382 -116 210 -72
rect 262 -65 1480 -64
rect 262 -116 1414 -65
rect -382 -117 1414 -116
rect 1466 -117 1480 -65
rect -382 -120 1480 -117
rect -382 -128 -370 -120
rect 203 -126 269 -120
rect 1407 -127 1473 -120
rect -450 -140 -370 -128
rect 30 -192 1980 -180
rect 30 -201 1912 -192
rect 30 -253 68 -201
rect 120 -253 478 -201
rect 530 -203 1277 -201
rect 530 -253 875 -203
rect 30 -255 875 -253
rect 927 -253 1277 -203
rect 1329 -248 1912 -201
rect 1968 -248 1980 -192
rect 1329 -253 1980 -248
rect 927 -255 1980 -253
rect 30 -260 1980 -255
rect 61 -263 127 -260
rect 471 -263 537 -260
rect 868 -265 934 -260
rect 1270 -263 1336 -260
rect 72 -2278 138 -2267
rect 72 -2280 79 -2278
rect -460 -2284 79 -2280
rect -460 -2336 -436 -2284
rect -384 -2330 79 -2284
rect 131 -2280 138 -2278
rect 1271 -2276 1337 -2265
rect 1271 -2280 1278 -2276
rect 131 -2328 1278 -2280
rect 1330 -2280 1337 -2276
rect 1330 -2328 1380 -2280
rect 131 -2330 1380 -2328
rect -384 -2336 1380 -2330
rect -460 -2340 1380 -2336
rect 475 -2400 541 -2392
rect 874 -2400 940 -2389
rect 2006 -2400 2072 -2392
rect -460 -2403 881 -2400
rect -460 -2455 482 -2403
rect 534 -2452 881 -2403
rect 933 -2403 2080 -2400
rect 933 -2452 2013 -2403
rect 534 -2455 2013 -2452
rect 2065 -2455 2080 -2403
rect -460 -2460 2080 -2455
rect 475 -2465 541 -2460
rect 874 -2462 940 -2460
rect 2006 -2465 2072 -2460
<< via2 >>
rect 1912 2312 1968 2368
rect 1092 2 1148 58
rect 1182 2 1238 58
rect -438 -128 -382 -72
rect 1912 -248 1968 -192
<< metal3 >>
rect 1900 2368 1980 2380
rect 1900 2312 1912 2368
rect 1968 2312 1980 2368
rect 1080 58 1250 70
rect 1080 2 1092 58
rect 1148 2 1182 58
rect 1238 2 1250 58
rect 1080 -10 1250 2
rect -450 -72 -370 -60
rect -450 -128 -438 -72
rect -382 -128 -370 -72
rect -450 -1750 -370 -128
rect -510 -1830 -370 -1750
rect 1130 -2970 1200 -10
rect 1900 -192 1980 2312
rect 1900 -248 1912 -192
rect 1968 -248 1980 -192
rect 1900 -260 1980 -248
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_0
timestamp 1757161594
transform 0 1 -252 -1 0 2544
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_1
timestamp 1757161594
transform 0 1 -252 -1 0 -2616
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_2
timestamp 1757161594
transform 0 1 148 -1 0 -2616
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_3
timestamp 1757161594
transform 0 1 548 -1 0 -2616
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_4
timestamp 1757161594
transform 0 1 948 -1 0 -2616
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_5
timestamp 1757161594
transform 0 1 1348 -1 0 -2616
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_6
timestamp 1757161594
transform 0 1 1748 -1 0 -2616
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_7
timestamp 1757161594
transform 0 1 1748 -1 0 2544
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_8
timestamp 1757161594
transform 0 1 1348 -1 0 2544
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_9
timestamp 1757161594
transform 0 1 948 -1 0 2544
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_10
timestamp 1757161594
transform 0 1 548 -1 0 2544
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_LHHU6U  sky130_fd_pr__pfet_01v8_lvt_LHHU6U_11
timestamp 1757161594
transform 0 1 148 -1 0 2544
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_0
timestamp 1757161594
transform 0 1 -252 -1 0 -1266
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_1
timestamp 1757161594
transform 0 1 148 -1 0 1294
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_2
timestamp 1757161594
transform 0 1 548 -1 0 1294
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_3
timestamp 1757161594
transform 0 1 948 -1 0 1294
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_4
timestamp 1757161594
transform 0 1 1348 -1 0 1294
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_5
timestamp 1757161594
transform 0 1 148 -1 0 -1266
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_6
timestamp 1757161594
transform 0 1 548 -1 0 -1266
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_7
timestamp 1757161594
transform 0 1 948 -1 0 -1266
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_8
timestamp 1757161594
transform 0 1 1348 -1 0 -1266
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_9
timestamp 1757161594
transform 0 1 1748 -1 0 -1266
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_10
timestamp 1757161594
transform 0 1 -252 -1 0 1294
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_W2HEQA  sky130_fd_pr__pfet_01v8_lvt_W2HEQA_11
timestamp 1757161594
transform 0 1 1748 -1 0 1294
box -1094 -148 1094 114
<< end >>
