magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< poly >>
rect -50 4414 50 4430
rect -50 4380 -17 4414
rect 17 4380 50 4414
rect -50 4000 50 4380
rect -50 -4380 50 -4000
rect -50 -4414 -17 -4380
rect 17 -4414 50 -4380
rect -50 -4430 50 -4414
<< polycont >>
rect -17 4380 17 4414
rect -17 -4414 17 -4380
<< npolyres >>
rect -50 -4000 50 4000
<< locali >>
rect -40 4380 -17 4414
rect 17 4380 40 4414
rect -34 4378 -17 4380
rect 17 4378 34 4380
rect -34 4340 34 4378
rect -34 4306 -17 4340
rect 17 4306 34 4340
rect -34 4268 34 4306
rect -34 4234 -17 4268
rect 17 4234 34 4268
rect -34 4196 34 4234
rect -34 4162 -17 4196
rect 17 4162 34 4196
rect -34 4124 34 4162
rect -34 4090 -17 4124
rect 17 4090 34 4124
rect -34 4052 34 4090
rect -34 4018 -17 4052
rect 17 4018 34 4052
rect -34 4017 34 4018
rect -34 -4019 34 -4017
rect -34 -4053 -17 -4019
rect 17 -4053 34 -4019
rect -34 -4091 34 -4053
rect -34 -4125 -17 -4091
rect 17 -4125 34 -4091
rect -34 -4163 34 -4125
rect -34 -4197 -17 -4163
rect 17 -4197 34 -4163
rect -34 -4235 34 -4197
rect -34 -4269 -17 -4235
rect 17 -4269 34 -4235
rect -34 -4307 34 -4269
rect -34 -4341 -17 -4307
rect 17 -4341 34 -4307
rect -34 -4379 34 -4341
rect -34 -4380 -17 -4379
rect 17 -4380 34 -4379
rect -40 -4414 -17 -4380
rect 17 -4414 40 -4380
<< viali >>
rect -17 4380 17 4412
rect -17 4378 17 4380
rect -17 4306 17 4340
rect -17 4234 17 4268
rect -17 4162 17 4196
rect -17 4090 17 4124
rect -17 4018 17 4052
rect -17 -4053 17 -4019
rect -17 -4125 17 -4091
rect -17 -4197 17 -4163
rect -17 -4269 17 -4235
rect -17 -4341 17 -4307
rect -17 -4380 17 -4379
rect -17 -4413 17 -4380
<< metal1 >>
rect -40 4412 40 4426
rect -40 4378 -17 4412
rect 17 4378 40 4412
rect -40 4340 40 4378
rect -40 4306 -17 4340
rect 17 4306 40 4340
rect -40 4268 40 4306
rect -40 4234 -17 4268
rect 17 4234 40 4268
rect -40 4196 40 4234
rect -40 4162 -17 4196
rect 17 4162 40 4196
rect -40 4124 40 4162
rect -40 4090 -17 4124
rect 17 4090 40 4124
rect -40 4052 40 4090
rect -40 4018 -17 4052
rect 17 4018 40 4052
rect -40 4005 40 4018
rect -40 -4019 40 -4005
rect -40 -4053 -17 -4019
rect 17 -4053 40 -4019
rect -40 -4091 40 -4053
rect -40 -4125 -17 -4091
rect 17 -4125 40 -4091
rect -40 -4163 40 -4125
rect -40 -4197 -17 -4163
rect 17 -4197 40 -4163
rect -40 -4235 40 -4197
rect -40 -4269 -17 -4235
rect 17 -4269 40 -4235
rect -40 -4307 40 -4269
rect -40 -4341 -17 -4307
rect 17 -4341 40 -4307
rect -40 -4379 40 -4341
rect -40 -4413 -17 -4379
rect 17 -4413 40 -4379
rect -40 -4426 40 -4413
<< end >>
