magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -184 -157 184 95
<< nmoslvt >>
rect -100 -131 100 69
<< ndiff >>
rect -158 20 -100 69
rect -158 -14 -146 20
rect -112 -14 -100 20
rect -158 -48 -100 -14
rect -158 -82 -146 -48
rect -112 -82 -100 -48
rect -158 -131 -100 -82
rect 100 20 158 69
rect 100 -14 112 20
rect 146 -14 158 20
rect 100 -48 158 -14
rect 100 -82 112 -48
rect 146 -82 158 -48
rect 100 -131 158 -82
<< ndiffc >>
rect -146 -14 -112 20
rect -146 -82 -112 -48
rect 112 -14 146 20
rect 112 -82 146 -48
<< poly >>
rect -75 141 75 157
rect -75 124 -51 141
rect -100 107 -51 124
rect -17 107 17 141
rect 51 124 75 141
rect 51 107 100 124
rect -100 69 100 107
rect -100 -157 100 -131
<< polycont >>
rect -51 107 -17 141
rect 17 107 51 141
<< locali >>
rect -75 107 -53 141
rect -17 107 17 141
rect 53 107 75 141
rect -146 22 -112 47
rect -146 -48 -112 -14
rect -146 -109 -112 -84
rect 112 22 146 47
rect 112 -48 146 -14
rect 112 -109 146 -84
<< viali >>
rect -53 107 -51 141
rect -51 107 -19 141
rect 19 107 51 141
rect 51 107 53 141
rect -146 20 -112 22
rect -146 -12 -112 20
rect -146 -82 -112 -50
rect -146 -84 -112 -82
rect 112 20 146 22
rect 112 -12 146 20
rect 112 -82 146 -50
rect 112 -84 146 -82
<< metal1 >>
rect -71 141 71 147
rect -71 107 -53 141
rect -19 107 19 141
rect 53 107 71 141
rect -71 101 71 107
rect -152 22 -106 43
rect -152 -12 -146 22
rect -112 -12 -106 22
rect -152 -50 -106 -12
rect -152 -84 -146 -50
rect -112 -84 -106 -50
rect -152 -105 -106 -84
rect 106 22 152 43
rect 106 -12 112 22
rect 146 -12 152 22
rect 106 -50 152 -12
rect 106 -84 112 -50
rect 146 -84 152 -50
rect 106 -105 152 -84
<< end >>
