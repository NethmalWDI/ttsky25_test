magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< error_s >>
rect -500 6738 -420 6750
rect -500 6682 -488 6738
rect -500 6670 -420 6682
rect -500 4478 -420 4490
rect -500 4422 -488 4478
rect -500 4410 -420 4422
<< pwell >>
rect -383 9287 3663 9373
rect -383 -507 -297 9287
rect 3577 -507 3663 9287
rect -383 -593 3663 -507
<< psubdiff >>
rect -357 9313 -281 9347
rect -247 9313 -213 9347
rect -179 9313 -145 9347
rect -111 9313 -77 9347
rect -43 9313 -9 9347
rect 25 9313 59 9347
rect 93 9313 127 9347
rect 161 9313 195 9347
rect 229 9313 263 9347
rect 297 9313 331 9347
rect 365 9313 399 9347
rect 433 9313 467 9347
rect 501 9313 535 9347
rect 569 9313 603 9347
rect 637 9313 671 9347
rect 705 9313 739 9347
rect 773 9313 807 9347
rect 841 9313 875 9347
rect 909 9313 943 9347
rect 977 9313 1011 9347
rect 1045 9313 1079 9347
rect 1113 9313 1147 9347
rect 1181 9313 1215 9347
rect 1249 9313 1283 9347
rect 1317 9313 1351 9347
rect 1385 9313 1419 9347
rect 1453 9313 1487 9347
rect 1521 9313 1555 9347
rect 1589 9313 1623 9347
rect 1657 9313 1691 9347
rect 1725 9313 1759 9347
rect 1793 9313 1827 9347
rect 1861 9313 1895 9347
rect 1929 9313 1963 9347
rect 1997 9313 2031 9347
rect 2065 9313 2099 9347
rect 2133 9313 2167 9347
rect 2201 9313 2235 9347
rect 2269 9313 2303 9347
rect 2337 9313 2371 9347
rect 2405 9313 2439 9347
rect 2473 9313 2507 9347
rect 2541 9313 2575 9347
rect 2609 9313 2643 9347
rect 2677 9313 2711 9347
rect 2745 9313 2779 9347
rect 2813 9313 2847 9347
rect 2881 9313 2915 9347
rect 2949 9313 2983 9347
rect 3017 9313 3051 9347
rect 3085 9313 3119 9347
rect 3153 9313 3187 9347
rect 3221 9313 3255 9347
rect 3289 9313 3323 9347
rect 3357 9313 3391 9347
rect 3425 9313 3459 9347
rect 3493 9313 3527 9347
rect 3561 9313 3637 9347
rect -357 9259 -323 9313
rect -357 9191 -323 9225
rect -357 9123 -323 9157
rect -357 9055 -323 9089
rect -357 8987 -323 9021
rect -357 8919 -323 8953
rect -357 8851 -323 8885
rect -357 8783 -323 8817
rect -357 8715 -323 8749
rect -357 8647 -323 8681
rect -357 8579 -323 8613
rect -357 8511 -323 8545
rect -357 8443 -323 8477
rect -357 8375 -323 8409
rect -357 8307 -323 8341
rect -357 8239 -323 8273
rect -357 8171 -323 8205
rect -357 8103 -323 8137
rect -357 8035 -323 8069
rect -357 7967 -323 8001
rect -357 7899 -323 7933
rect -357 7831 -323 7865
rect -357 7763 -323 7797
rect -357 7695 -323 7729
rect -357 7627 -323 7661
rect -357 7559 -323 7593
rect -357 7491 -323 7525
rect -357 7423 -323 7457
rect -357 7355 -323 7389
rect -357 7287 -323 7321
rect -357 7219 -323 7253
rect -357 7151 -323 7185
rect -357 7083 -323 7117
rect -357 7015 -323 7049
rect -357 6947 -323 6981
rect -357 6879 -323 6913
rect -357 6811 -323 6845
rect -357 6743 -323 6777
rect -357 6675 -323 6709
rect -357 6607 -323 6641
rect -357 6539 -323 6573
rect -357 6471 -323 6505
rect -357 6403 -323 6437
rect -357 6335 -323 6369
rect -357 6267 -323 6301
rect -357 6199 -323 6233
rect -357 6131 -323 6165
rect -357 6063 -323 6097
rect -357 5995 -323 6029
rect -357 5927 -323 5961
rect -357 5859 -323 5893
rect -357 5791 -323 5825
rect -357 5723 -323 5757
rect -357 5655 -323 5689
rect -357 5587 -323 5621
rect -357 5519 -323 5553
rect -357 5451 -323 5485
rect -357 5383 -323 5417
rect -357 5315 -323 5349
rect -357 5247 -323 5281
rect -357 5179 -323 5213
rect -357 5111 -323 5145
rect -357 5043 -323 5077
rect -357 4975 -323 5009
rect -357 4907 -323 4941
rect -357 4839 -323 4873
rect -357 4771 -323 4805
rect -357 4703 -323 4737
rect -357 4635 -323 4669
rect -357 4567 -323 4601
rect -357 4499 -323 4533
rect -357 4431 -323 4465
rect -357 4363 -323 4397
rect -357 4295 -323 4329
rect -357 4227 -323 4261
rect -357 4159 -323 4193
rect -357 4091 -323 4125
rect -357 4023 -323 4057
rect -357 3955 -323 3989
rect -357 3887 -323 3921
rect -357 3819 -323 3853
rect -357 3751 -323 3785
rect -357 3683 -323 3717
rect -357 3615 -323 3649
rect -357 3547 -323 3581
rect -357 3479 -323 3513
rect -357 3411 -323 3445
rect -357 3343 -323 3377
rect -357 3275 -323 3309
rect -357 3207 -323 3241
rect -357 3139 -323 3173
rect -357 3071 -323 3105
rect -357 3003 -323 3037
rect -357 2935 -323 2969
rect -357 2867 -323 2901
rect -357 2799 -323 2833
rect -357 2731 -323 2765
rect -357 2663 -323 2697
rect -357 2595 -323 2629
rect -357 2527 -323 2561
rect -357 2459 -323 2493
rect -357 2391 -323 2425
rect -357 2323 -323 2357
rect -357 2255 -323 2289
rect -357 2187 -323 2221
rect -357 2119 -323 2153
rect -357 2051 -323 2085
rect -357 1983 -323 2017
rect -357 1915 -323 1949
rect -357 1847 -323 1881
rect -357 1779 -323 1813
rect -357 1711 -323 1745
rect -357 1643 -323 1677
rect -357 1575 -323 1609
rect -357 1507 -323 1541
rect -357 1439 -323 1473
rect -357 1371 -323 1405
rect -357 1303 -323 1337
rect -357 1235 -323 1269
rect -357 1167 -323 1201
rect -357 1099 -323 1133
rect -357 1031 -323 1065
rect -357 963 -323 997
rect -357 895 -323 929
rect -357 827 -323 861
rect -357 759 -323 793
rect -357 691 -323 725
rect -357 623 -323 657
rect -357 555 -323 589
rect -357 487 -323 521
rect -357 419 -323 453
rect -357 351 -323 385
rect -357 283 -323 317
rect -357 215 -323 249
rect -357 147 -323 181
rect -357 79 -323 113
rect -357 11 -323 45
rect -357 -57 -323 -23
rect -357 -125 -323 -91
rect -357 -193 -323 -159
rect -357 -261 -323 -227
rect -357 -329 -323 -295
rect -357 -397 -323 -363
rect -357 -465 -323 -431
rect -357 -533 -323 -499
rect 3603 9259 3637 9313
rect 3603 9191 3637 9225
rect 3603 9123 3637 9157
rect 3603 9055 3637 9089
rect 3603 8987 3637 9021
rect 3603 8919 3637 8953
rect 3603 8851 3637 8885
rect 3603 8783 3637 8817
rect 3603 8715 3637 8749
rect 3603 8647 3637 8681
rect 3603 8579 3637 8613
rect 3603 8511 3637 8545
rect 3603 8443 3637 8477
rect 3603 8375 3637 8409
rect 3603 8307 3637 8341
rect 3603 8239 3637 8273
rect 3603 8171 3637 8205
rect 3603 8103 3637 8137
rect 3603 8035 3637 8069
rect 3603 7967 3637 8001
rect 3603 7899 3637 7933
rect 3603 7831 3637 7865
rect 3603 7763 3637 7797
rect 3603 7695 3637 7729
rect 3603 7627 3637 7661
rect 3603 7559 3637 7593
rect 3603 7491 3637 7525
rect 3603 7423 3637 7457
rect 3603 7355 3637 7389
rect 3603 7287 3637 7321
rect 3603 7219 3637 7253
rect 3603 7151 3637 7185
rect 3603 7083 3637 7117
rect 3603 7015 3637 7049
rect 3603 6947 3637 6981
rect 3603 6879 3637 6913
rect 3603 6811 3637 6845
rect 3603 6743 3637 6777
rect 3603 6675 3637 6709
rect 3603 6607 3637 6641
rect 3603 6539 3637 6573
rect 3603 6471 3637 6505
rect 3603 6403 3637 6437
rect 3603 6335 3637 6369
rect 3603 6267 3637 6301
rect 3603 6199 3637 6233
rect 3603 6131 3637 6165
rect 3603 6063 3637 6097
rect 3603 5995 3637 6029
rect 3603 5927 3637 5961
rect 3603 5859 3637 5893
rect 3603 5791 3637 5825
rect 3603 5723 3637 5757
rect 3603 5655 3637 5689
rect 3603 5587 3637 5621
rect 3603 5519 3637 5553
rect 3603 5451 3637 5485
rect 3603 5383 3637 5417
rect 3603 5315 3637 5349
rect 3603 5247 3637 5281
rect 3603 5179 3637 5213
rect 3603 5111 3637 5145
rect 3603 5043 3637 5077
rect 3603 4975 3637 5009
rect 3603 4907 3637 4941
rect 3603 4839 3637 4873
rect 3603 4771 3637 4805
rect 3603 4703 3637 4737
rect 3603 4635 3637 4669
rect 3603 4567 3637 4601
rect 3603 4499 3637 4533
rect 3603 4431 3637 4465
rect 3603 4363 3637 4397
rect 3603 4295 3637 4329
rect 3603 4227 3637 4261
rect 3603 4159 3637 4193
rect 3603 4091 3637 4125
rect 3603 4023 3637 4057
rect 3603 3955 3637 3989
rect 3603 3887 3637 3921
rect 3603 3819 3637 3853
rect 3603 3751 3637 3785
rect 3603 3683 3637 3717
rect 3603 3615 3637 3649
rect 3603 3547 3637 3581
rect 3603 3479 3637 3513
rect 3603 3411 3637 3445
rect 3603 3343 3637 3377
rect 3603 3275 3637 3309
rect 3603 3207 3637 3241
rect 3603 3139 3637 3173
rect 3603 3071 3637 3105
rect 3603 3003 3637 3037
rect 3603 2935 3637 2969
rect 3603 2867 3637 2901
rect 3603 2799 3637 2833
rect 3603 2731 3637 2765
rect 3603 2663 3637 2697
rect 3603 2595 3637 2629
rect 3603 2527 3637 2561
rect 3603 2459 3637 2493
rect 3603 2391 3637 2425
rect 3603 2323 3637 2357
rect 3603 2255 3637 2289
rect 3603 2187 3637 2221
rect 3603 2119 3637 2153
rect 3603 2051 3637 2085
rect 3603 1983 3637 2017
rect 3603 1915 3637 1949
rect 3603 1847 3637 1881
rect 3603 1779 3637 1813
rect 3603 1711 3637 1745
rect 3603 1643 3637 1677
rect 3603 1575 3637 1609
rect 3603 1507 3637 1541
rect 3603 1439 3637 1473
rect 3603 1371 3637 1405
rect 3603 1303 3637 1337
rect 3603 1235 3637 1269
rect 3603 1167 3637 1201
rect 3603 1099 3637 1133
rect 3603 1031 3637 1065
rect 3603 963 3637 997
rect 3603 895 3637 929
rect 3603 827 3637 861
rect 3603 759 3637 793
rect 3603 691 3637 725
rect 3603 623 3637 657
rect 3603 555 3637 589
rect 3603 487 3637 521
rect 3603 419 3637 453
rect 3603 351 3637 385
rect 3603 283 3637 317
rect 3603 215 3637 249
rect 3603 147 3637 181
rect 3603 79 3637 113
rect 3603 11 3637 45
rect 3603 -57 3637 -23
rect 3603 -125 3637 -91
rect 3603 -193 3637 -159
rect 3603 -261 3637 -227
rect 3603 -329 3637 -295
rect 3603 -397 3637 -363
rect 3603 -465 3637 -431
rect 3603 -533 3637 -499
rect -357 -567 -281 -533
rect -247 -567 -213 -533
rect -179 -567 -145 -533
rect -111 -567 -77 -533
rect -43 -567 -9 -533
rect 25 -567 59 -533
rect 93 -567 127 -533
rect 161 -567 195 -533
rect 229 -567 263 -533
rect 297 -567 331 -533
rect 365 -567 399 -533
rect 433 -567 467 -533
rect 501 -567 535 -533
rect 569 -567 603 -533
rect 637 -567 671 -533
rect 705 -567 739 -533
rect 773 -567 807 -533
rect 841 -567 875 -533
rect 909 -567 943 -533
rect 977 -567 1011 -533
rect 1045 -567 1079 -533
rect 1113 -567 1147 -533
rect 1181 -567 1215 -533
rect 1249 -567 1283 -533
rect 1317 -567 1351 -533
rect 1385 -567 1419 -533
rect 1453 -567 1487 -533
rect 1521 -567 1555 -533
rect 1589 -567 1623 -533
rect 1657 -567 1691 -533
rect 1725 -567 1759 -533
rect 1793 -567 1827 -533
rect 1861 -567 1895 -533
rect 1929 -567 1963 -533
rect 1997 -567 2031 -533
rect 2065 -567 2099 -533
rect 2133 -567 2167 -533
rect 2201 -567 2235 -533
rect 2269 -567 2303 -533
rect 2337 -567 2371 -533
rect 2405 -567 2439 -533
rect 2473 -567 2507 -533
rect 2541 -567 2575 -533
rect 2609 -567 2643 -533
rect 2677 -567 2711 -533
rect 2745 -567 2779 -533
rect 2813 -567 2847 -533
rect 2881 -567 2915 -533
rect 2949 -567 2983 -533
rect 3017 -567 3051 -533
rect 3085 -567 3119 -533
rect 3153 -567 3187 -533
rect 3221 -567 3255 -533
rect 3289 -567 3323 -533
rect 3357 -567 3391 -533
rect 3425 -567 3459 -533
rect 3493 -567 3527 -533
rect 3561 -567 3637 -533
<< psubdiffcont >>
rect -281 9313 -247 9347
rect -213 9313 -179 9347
rect -145 9313 -111 9347
rect -77 9313 -43 9347
rect -9 9313 25 9347
rect 59 9313 93 9347
rect 127 9313 161 9347
rect 195 9313 229 9347
rect 263 9313 297 9347
rect 331 9313 365 9347
rect 399 9313 433 9347
rect 467 9313 501 9347
rect 535 9313 569 9347
rect 603 9313 637 9347
rect 671 9313 705 9347
rect 739 9313 773 9347
rect 807 9313 841 9347
rect 875 9313 909 9347
rect 943 9313 977 9347
rect 1011 9313 1045 9347
rect 1079 9313 1113 9347
rect 1147 9313 1181 9347
rect 1215 9313 1249 9347
rect 1283 9313 1317 9347
rect 1351 9313 1385 9347
rect 1419 9313 1453 9347
rect 1487 9313 1521 9347
rect 1555 9313 1589 9347
rect 1623 9313 1657 9347
rect 1691 9313 1725 9347
rect 1759 9313 1793 9347
rect 1827 9313 1861 9347
rect 1895 9313 1929 9347
rect 1963 9313 1997 9347
rect 2031 9313 2065 9347
rect 2099 9313 2133 9347
rect 2167 9313 2201 9347
rect 2235 9313 2269 9347
rect 2303 9313 2337 9347
rect 2371 9313 2405 9347
rect 2439 9313 2473 9347
rect 2507 9313 2541 9347
rect 2575 9313 2609 9347
rect 2643 9313 2677 9347
rect 2711 9313 2745 9347
rect 2779 9313 2813 9347
rect 2847 9313 2881 9347
rect 2915 9313 2949 9347
rect 2983 9313 3017 9347
rect 3051 9313 3085 9347
rect 3119 9313 3153 9347
rect 3187 9313 3221 9347
rect 3255 9313 3289 9347
rect 3323 9313 3357 9347
rect 3391 9313 3425 9347
rect 3459 9313 3493 9347
rect 3527 9313 3561 9347
rect -357 9225 -323 9259
rect -357 9157 -323 9191
rect -357 9089 -323 9123
rect -357 9021 -323 9055
rect -357 8953 -323 8987
rect -357 8885 -323 8919
rect -357 8817 -323 8851
rect -357 8749 -323 8783
rect -357 8681 -323 8715
rect -357 8613 -323 8647
rect -357 8545 -323 8579
rect -357 8477 -323 8511
rect -357 8409 -323 8443
rect -357 8341 -323 8375
rect -357 8273 -323 8307
rect -357 8205 -323 8239
rect -357 8137 -323 8171
rect -357 8069 -323 8103
rect -357 8001 -323 8035
rect -357 7933 -323 7967
rect -357 7865 -323 7899
rect -357 7797 -323 7831
rect -357 7729 -323 7763
rect -357 7661 -323 7695
rect -357 7593 -323 7627
rect -357 7525 -323 7559
rect -357 7457 -323 7491
rect -357 7389 -323 7423
rect -357 7321 -323 7355
rect -357 7253 -323 7287
rect -357 7185 -323 7219
rect -357 7117 -323 7151
rect -357 7049 -323 7083
rect -357 6981 -323 7015
rect -357 6913 -323 6947
rect -357 6845 -323 6879
rect -357 6777 -323 6811
rect -357 6709 -323 6743
rect -357 6641 -323 6675
rect -357 6573 -323 6607
rect -357 6505 -323 6539
rect -357 6437 -323 6471
rect -357 6369 -323 6403
rect -357 6301 -323 6335
rect -357 6233 -323 6267
rect -357 6165 -323 6199
rect -357 6097 -323 6131
rect -357 6029 -323 6063
rect -357 5961 -323 5995
rect -357 5893 -323 5927
rect -357 5825 -323 5859
rect -357 5757 -323 5791
rect -357 5689 -323 5723
rect -357 5621 -323 5655
rect -357 5553 -323 5587
rect -357 5485 -323 5519
rect -357 5417 -323 5451
rect -357 5349 -323 5383
rect -357 5281 -323 5315
rect -357 5213 -323 5247
rect -357 5145 -323 5179
rect -357 5077 -323 5111
rect -357 5009 -323 5043
rect -357 4941 -323 4975
rect -357 4873 -323 4907
rect -357 4805 -323 4839
rect -357 4737 -323 4771
rect -357 4669 -323 4703
rect -357 4601 -323 4635
rect -357 4533 -323 4567
rect -357 4465 -323 4499
rect -357 4397 -323 4431
rect -357 4329 -323 4363
rect -357 4261 -323 4295
rect -357 4193 -323 4227
rect -357 4125 -323 4159
rect -357 4057 -323 4091
rect -357 3989 -323 4023
rect -357 3921 -323 3955
rect -357 3853 -323 3887
rect -357 3785 -323 3819
rect -357 3717 -323 3751
rect -357 3649 -323 3683
rect -357 3581 -323 3615
rect -357 3513 -323 3547
rect -357 3445 -323 3479
rect -357 3377 -323 3411
rect -357 3309 -323 3343
rect -357 3241 -323 3275
rect -357 3173 -323 3207
rect -357 3105 -323 3139
rect -357 3037 -323 3071
rect -357 2969 -323 3003
rect -357 2901 -323 2935
rect -357 2833 -323 2867
rect -357 2765 -323 2799
rect -357 2697 -323 2731
rect -357 2629 -323 2663
rect -357 2561 -323 2595
rect -357 2493 -323 2527
rect -357 2425 -323 2459
rect -357 2357 -323 2391
rect -357 2289 -323 2323
rect -357 2221 -323 2255
rect -357 2153 -323 2187
rect -357 2085 -323 2119
rect -357 2017 -323 2051
rect -357 1949 -323 1983
rect -357 1881 -323 1915
rect -357 1813 -323 1847
rect -357 1745 -323 1779
rect -357 1677 -323 1711
rect -357 1609 -323 1643
rect -357 1541 -323 1575
rect -357 1473 -323 1507
rect -357 1405 -323 1439
rect -357 1337 -323 1371
rect -357 1269 -323 1303
rect -357 1201 -323 1235
rect -357 1133 -323 1167
rect -357 1065 -323 1099
rect -357 997 -323 1031
rect -357 929 -323 963
rect -357 861 -323 895
rect -357 793 -323 827
rect -357 725 -323 759
rect -357 657 -323 691
rect -357 589 -323 623
rect -357 521 -323 555
rect -357 453 -323 487
rect -357 385 -323 419
rect -357 317 -323 351
rect -357 249 -323 283
rect -357 181 -323 215
rect -357 113 -323 147
rect -357 45 -323 79
rect -357 -23 -323 11
rect -357 -91 -323 -57
rect -357 -159 -323 -125
rect -357 -227 -323 -193
rect -357 -295 -323 -261
rect -357 -363 -323 -329
rect -357 -431 -323 -397
rect -357 -499 -323 -465
rect 3603 9225 3637 9259
rect 3603 9157 3637 9191
rect 3603 9089 3637 9123
rect 3603 9021 3637 9055
rect 3603 8953 3637 8987
rect 3603 8885 3637 8919
rect 3603 8817 3637 8851
rect 3603 8749 3637 8783
rect 3603 8681 3637 8715
rect 3603 8613 3637 8647
rect 3603 8545 3637 8579
rect 3603 8477 3637 8511
rect 3603 8409 3637 8443
rect 3603 8341 3637 8375
rect 3603 8273 3637 8307
rect 3603 8205 3637 8239
rect 3603 8137 3637 8171
rect 3603 8069 3637 8103
rect 3603 8001 3637 8035
rect 3603 7933 3637 7967
rect 3603 7865 3637 7899
rect 3603 7797 3637 7831
rect 3603 7729 3637 7763
rect 3603 7661 3637 7695
rect 3603 7593 3637 7627
rect 3603 7525 3637 7559
rect 3603 7457 3637 7491
rect 3603 7389 3637 7423
rect 3603 7321 3637 7355
rect 3603 7253 3637 7287
rect 3603 7185 3637 7219
rect 3603 7117 3637 7151
rect 3603 7049 3637 7083
rect 3603 6981 3637 7015
rect 3603 6913 3637 6947
rect 3603 6845 3637 6879
rect 3603 6777 3637 6811
rect 3603 6709 3637 6743
rect 3603 6641 3637 6675
rect 3603 6573 3637 6607
rect 3603 6505 3637 6539
rect 3603 6437 3637 6471
rect 3603 6369 3637 6403
rect 3603 6301 3637 6335
rect 3603 6233 3637 6267
rect 3603 6165 3637 6199
rect 3603 6097 3637 6131
rect 3603 6029 3637 6063
rect 3603 5961 3637 5995
rect 3603 5893 3637 5927
rect 3603 5825 3637 5859
rect 3603 5757 3637 5791
rect 3603 5689 3637 5723
rect 3603 5621 3637 5655
rect 3603 5553 3637 5587
rect 3603 5485 3637 5519
rect 3603 5417 3637 5451
rect 3603 5349 3637 5383
rect 3603 5281 3637 5315
rect 3603 5213 3637 5247
rect 3603 5145 3637 5179
rect 3603 5077 3637 5111
rect 3603 5009 3637 5043
rect 3603 4941 3637 4975
rect 3603 4873 3637 4907
rect 3603 4805 3637 4839
rect 3603 4737 3637 4771
rect 3603 4669 3637 4703
rect 3603 4601 3637 4635
rect 3603 4533 3637 4567
rect 3603 4465 3637 4499
rect 3603 4397 3637 4431
rect 3603 4329 3637 4363
rect 3603 4261 3637 4295
rect 3603 4193 3637 4227
rect 3603 4125 3637 4159
rect 3603 4057 3637 4091
rect 3603 3989 3637 4023
rect 3603 3921 3637 3955
rect 3603 3853 3637 3887
rect 3603 3785 3637 3819
rect 3603 3717 3637 3751
rect 3603 3649 3637 3683
rect 3603 3581 3637 3615
rect 3603 3513 3637 3547
rect 3603 3445 3637 3479
rect 3603 3377 3637 3411
rect 3603 3309 3637 3343
rect 3603 3241 3637 3275
rect 3603 3173 3637 3207
rect 3603 3105 3637 3139
rect 3603 3037 3637 3071
rect 3603 2969 3637 3003
rect 3603 2901 3637 2935
rect 3603 2833 3637 2867
rect 3603 2765 3637 2799
rect 3603 2697 3637 2731
rect 3603 2629 3637 2663
rect 3603 2561 3637 2595
rect 3603 2493 3637 2527
rect 3603 2425 3637 2459
rect 3603 2357 3637 2391
rect 3603 2289 3637 2323
rect 3603 2221 3637 2255
rect 3603 2153 3637 2187
rect 3603 2085 3637 2119
rect 3603 2017 3637 2051
rect 3603 1949 3637 1983
rect 3603 1881 3637 1915
rect 3603 1813 3637 1847
rect 3603 1745 3637 1779
rect 3603 1677 3637 1711
rect 3603 1609 3637 1643
rect 3603 1541 3637 1575
rect 3603 1473 3637 1507
rect 3603 1405 3637 1439
rect 3603 1337 3637 1371
rect 3603 1269 3637 1303
rect 3603 1201 3637 1235
rect 3603 1133 3637 1167
rect 3603 1065 3637 1099
rect 3603 997 3637 1031
rect 3603 929 3637 963
rect 3603 861 3637 895
rect 3603 793 3637 827
rect 3603 725 3637 759
rect 3603 657 3637 691
rect 3603 589 3637 623
rect 3603 521 3637 555
rect 3603 453 3637 487
rect 3603 385 3637 419
rect 3603 317 3637 351
rect 3603 249 3637 283
rect 3603 181 3637 215
rect 3603 113 3637 147
rect 3603 45 3637 79
rect 3603 -23 3637 11
rect 3603 -91 3637 -57
rect 3603 -159 3637 -125
rect 3603 -227 3637 -193
rect 3603 -295 3637 -261
rect 3603 -363 3637 -329
rect 3603 -431 3637 -397
rect 3603 -499 3637 -465
rect -281 -567 -247 -533
rect -213 -567 -179 -533
rect -145 -567 -111 -533
rect -77 -567 -43 -533
rect -9 -567 25 -533
rect 59 -567 93 -533
rect 127 -567 161 -533
rect 195 -567 229 -533
rect 263 -567 297 -533
rect 331 -567 365 -533
rect 399 -567 433 -533
rect 467 -567 501 -533
rect 535 -567 569 -533
rect 603 -567 637 -533
rect 671 -567 705 -533
rect 739 -567 773 -533
rect 807 -567 841 -533
rect 875 -567 909 -533
rect 943 -567 977 -533
rect 1011 -567 1045 -533
rect 1079 -567 1113 -533
rect 1147 -567 1181 -533
rect 1215 -567 1249 -533
rect 1283 -567 1317 -533
rect 1351 -567 1385 -533
rect 1419 -567 1453 -533
rect 1487 -567 1521 -533
rect 1555 -567 1589 -533
rect 1623 -567 1657 -533
rect 1691 -567 1725 -533
rect 1759 -567 1793 -533
rect 1827 -567 1861 -533
rect 1895 -567 1929 -533
rect 1963 -567 1997 -533
rect 2031 -567 2065 -533
rect 2099 -567 2133 -533
rect 2167 -567 2201 -533
rect 2235 -567 2269 -533
rect 2303 -567 2337 -533
rect 2371 -567 2405 -533
rect 2439 -567 2473 -533
rect 2507 -567 2541 -533
rect 2575 -567 2609 -533
rect 2643 -567 2677 -533
rect 2711 -567 2745 -533
rect 2779 -567 2813 -533
rect 2847 -567 2881 -533
rect 2915 -567 2949 -533
rect 2983 -567 3017 -533
rect 3051 -567 3085 -533
rect 3119 -567 3153 -533
rect 3187 -567 3221 -533
rect 3255 -567 3289 -533
rect 3323 -567 3357 -533
rect 3391 -567 3425 -533
rect 3459 -567 3493 -533
rect 3527 -567 3561 -533
<< locali >>
rect -357 9313 -281 9347
rect -247 9313 -213 9347
rect -179 9313 -145 9347
rect -111 9313 -77 9347
rect -43 9313 -9 9347
rect 25 9313 59 9347
rect 93 9313 127 9347
rect 161 9313 195 9347
rect 229 9313 263 9347
rect 297 9313 331 9347
rect 365 9313 399 9347
rect 433 9313 467 9347
rect 501 9313 535 9347
rect 569 9313 603 9347
rect 637 9313 671 9347
rect 705 9313 739 9347
rect 773 9313 807 9347
rect 841 9313 875 9347
rect 909 9313 943 9347
rect 977 9313 1011 9347
rect 1045 9313 1079 9347
rect 1113 9313 1147 9347
rect 1181 9313 1215 9347
rect 1249 9313 1283 9347
rect 1317 9313 1351 9347
rect 1385 9313 1419 9347
rect 1453 9313 1487 9347
rect 1521 9313 1555 9347
rect 1589 9313 1623 9347
rect 1657 9313 1691 9347
rect 1725 9313 1759 9347
rect 1793 9313 1827 9347
rect 1861 9313 1895 9347
rect 1929 9313 1963 9347
rect 1997 9313 2031 9347
rect 2065 9313 2099 9347
rect 2133 9313 2167 9347
rect 2201 9313 2235 9347
rect 2269 9313 2303 9347
rect 2337 9313 2371 9347
rect 2405 9313 2439 9347
rect 2473 9313 2507 9347
rect 2541 9313 2575 9347
rect 2609 9313 2643 9347
rect 2677 9313 2711 9347
rect 2745 9313 2779 9347
rect 2813 9313 2847 9347
rect 2881 9313 2915 9347
rect 2949 9313 2983 9347
rect 3017 9313 3051 9347
rect 3085 9313 3119 9347
rect 3153 9313 3187 9347
rect 3221 9313 3255 9347
rect 3289 9313 3323 9347
rect 3357 9313 3391 9347
rect 3425 9313 3459 9347
rect 3493 9313 3527 9347
rect 3561 9313 3637 9347
rect -357 9259 -323 9313
rect -357 9191 -323 9225
rect -357 9123 -323 9157
rect -357 9055 -323 9089
rect -357 8987 -323 9021
rect -357 8919 -323 8953
rect -357 8851 -323 8885
rect -357 8783 -323 8817
rect -357 8715 -323 8749
rect -357 8647 -323 8681
rect -357 8579 -323 8613
rect -357 8511 -323 8545
rect -357 8443 -323 8477
rect -357 8375 -323 8409
rect -357 8307 -323 8341
rect -357 8239 -323 8273
rect -357 8171 -323 8205
rect -357 8103 -323 8137
rect -357 8035 -323 8069
rect -357 7967 -323 8001
rect -357 7899 -323 7933
rect -357 7831 -323 7865
rect -357 7763 -323 7797
rect -357 7695 -323 7729
rect -357 7627 -323 7661
rect -357 7559 -323 7593
rect -357 7491 -323 7525
rect -357 7423 -323 7457
rect -357 7355 -323 7389
rect -357 7287 -323 7321
rect -357 7219 -323 7253
rect -357 7151 -323 7185
rect -357 7083 -323 7117
rect -357 7015 -323 7049
rect -357 6947 -323 6981
rect -357 6879 -323 6913
rect -357 6811 -323 6845
rect -357 6743 -323 6777
rect -357 6675 -323 6709
rect -357 6607 -323 6641
rect -357 6539 -323 6573
rect -357 6471 -323 6505
rect -357 6403 -323 6437
rect -357 6335 -323 6369
rect -357 6267 -323 6301
rect -357 6199 -323 6233
rect -357 6131 -323 6165
rect -357 6063 -323 6097
rect -357 5995 -323 6029
rect -357 5927 -323 5961
rect -357 5859 -323 5893
rect -357 5791 -323 5825
rect -357 5723 -323 5757
rect -357 5655 -323 5689
rect -357 5587 -323 5621
rect -357 5519 -323 5553
rect -357 5451 -323 5485
rect -357 5383 -323 5417
rect -357 5315 -323 5349
rect -357 5247 -323 5281
rect -357 5179 -323 5213
rect -357 5111 -323 5145
rect -357 5043 -323 5077
rect -357 4975 -323 5009
rect -357 4907 -323 4941
rect -357 4839 -323 4873
rect -357 4771 -323 4805
rect -357 4703 -323 4737
rect -357 4635 -323 4669
rect -357 4567 -323 4601
rect -357 4499 -323 4533
rect -357 4431 -323 4465
rect -357 4363 -323 4397
rect -357 4295 -323 4329
rect -357 4227 -323 4261
rect -357 4159 -323 4193
rect -357 4091 -323 4125
rect -357 4023 -323 4057
rect -357 3955 -323 3989
rect -357 3887 -323 3921
rect -357 3819 -323 3853
rect -357 3751 -323 3785
rect -357 3683 -323 3717
rect -357 3615 -323 3649
rect -357 3547 -323 3581
rect -357 3479 -323 3513
rect -357 3411 -323 3445
rect -357 3343 -323 3377
rect -357 3275 -323 3309
rect -357 3207 -323 3241
rect -357 3139 -323 3173
rect -357 3071 -323 3105
rect -357 3003 -323 3037
rect -357 2935 -323 2969
rect -357 2867 -323 2901
rect -357 2799 -323 2833
rect -357 2731 -323 2765
rect -357 2663 -323 2697
rect -357 2595 -323 2629
rect -357 2527 -323 2561
rect -357 2459 -323 2493
rect -357 2391 -323 2425
rect -357 2323 -323 2357
rect -357 2255 -323 2289
rect -357 2187 -323 2221
rect -357 2119 -323 2153
rect -357 2051 -323 2085
rect -357 1983 -323 2017
rect -357 1915 -323 1949
rect -357 1847 -323 1881
rect -357 1779 -323 1813
rect -357 1711 -323 1745
rect -357 1643 -323 1677
rect -357 1575 -323 1609
rect -357 1507 -323 1541
rect -357 1439 -323 1473
rect -357 1371 -323 1405
rect -357 1303 -323 1337
rect -357 1235 -323 1269
rect -357 1167 -323 1201
rect -357 1099 -323 1133
rect -357 1031 -323 1065
rect -357 963 -323 997
rect -357 895 -323 929
rect -357 827 -323 861
rect -357 759 -323 793
rect -357 691 -323 725
rect -357 623 -323 657
rect -357 555 -323 589
rect -357 487 -323 521
rect -357 419 -323 453
rect -357 351 -323 385
rect -357 283 -323 317
rect -357 215 -323 249
rect -357 147 -323 181
rect -357 79 -323 113
rect -357 11 -323 45
rect -357 -57 -323 -23
rect -357 -125 -323 -91
rect -357 -193 -323 -159
rect -357 -261 -323 -227
rect -357 -329 -323 -295
rect -357 -397 -323 -363
rect -357 -465 -323 -431
rect -357 -533 -323 -499
rect 3603 9259 3637 9313
rect 3603 9191 3637 9225
rect 3603 9123 3637 9157
rect 3603 9055 3637 9089
rect 3603 8987 3637 9021
rect 3603 8919 3637 8953
rect 3603 8851 3637 8885
rect 3603 8783 3637 8817
rect 3603 8715 3637 8749
rect 3603 8647 3637 8681
rect 3603 8579 3637 8613
rect 3603 8511 3637 8545
rect 3603 8443 3637 8477
rect 3603 8375 3637 8409
rect 3603 8307 3637 8341
rect 3603 8239 3637 8273
rect 3603 8171 3637 8205
rect 3603 8103 3637 8137
rect 3603 8035 3637 8069
rect 3603 7967 3637 8001
rect 3603 7899 3637 7933
rect 3603 7831 3637 7865
rect 3603 7763 3637 7797
rect 3603 7695 3637 7729
rect 3603 7627 3637 7661
rect 3603 7559 3637 7593
rect 3603 7491 3637 7525
rect 3603 7423 3637 7457
rect 3603 7355 3637 7389
rect 3603 7287 3637 7321
rect 3603 7219 3637 7253
rect 3603 7151 3637 7185
rect 3603 7083 3637 7117
rect 3603 7015 3637 7049
rect 3603 6947 3637 6981
rect 3603 6879 3637 6913
rect 3603 6811 3637 6845
rect 3603 6743 3637 6777
rect 3603 6675 3637 6709
rect 3603 6607 3637 6641
rect 3603 6539 3637 6573
rect 3603 6471 3637 6505
rect 3603 6403 3637 6437
rect 3603 6335 3637 6369
rect 3603 6267 3637 6301
rect 3603 6199 3637 6233
rect 3603 6131 3637 6165
rect 3603 6063 3637 6097
rect 3603 5995 3637 6029
rect 3603 5927 3637 5961
rect 3603 5859 3637 5893
rect 3603 5791 3637 5825
rect 3603 5723 3637 5757
rect 3603 5655 3637 5689
rect 3603 5587 3637 5621
rect 3603 5519 3637 5553
rect 3603 5451 3637 5485
rect 3603 5383 3637 5417
rect 3603 5315 3637 5349
rect 3603 5247 3637 5281
rect 3603 5179 3637 5213
rect 3603 5111 3637 5145
rect 3603 5043 3637 5077
rect 3603 4975 3637 5009
rect 3603 4907 3637 4941
rect 3603 4839 3637 4873
rect 3603 4771 3637 4805
rect 3603 4703 3637 4737
rect 3603 4635 3637 4669
rect 3603 4567 3637 4601
rect 3603 4499 3637 4533
rect 3603 4431 3637 4465
rect 3603 4363 3637 4397
rect 3603 4295 3637 4329
rect 3603 4227 3637 4261
rect 3603 4159 3637 4193
rect 3603 4091 3637 4125
rect 3603 4023 3637 4057
rect 3603 3955 3637 3989
rect 3603 3887 3637 3921
rect 3603 3819 3637 3853
rect 3603 3751 3637 3785
rect 3603 3683 3637 3717
rect 3603 3615 3637 3649
rect 3603 3547 3637 3581
rect 3603 3479 3637 3513
rect 3603 3411 3637 3445
rect 3603 3343 3637 3377
rect 3603 3275 3637 3309
rect 3603 3207 3637 3241
rect 3603 3139 3637 3173
rect 3603 3071 3637 3105
rect 3603 3003 3637 3037
rect 3603 2935 3637 2969
rect 3603 2867 3637 2901
rect 3603 2799 3637 2833
rect 3603 2731 3637 2765
rect 3603 2663 3637 2697
rect 3603 2595 3637 2629
rect 3603 2527 3637 2561
rect 3603 2459 3637 2493
rect 3603 2391 3637 2425
rect 3603 2323 3637 2357
rect 3603 2255 3637 2289
rect 3603 2187 3637 2221
rect 3603 2119 3637 2153
rect 3603 2051 3637 2085
rect 3603 1983 3637 2017
rect 3603 1915 3637 1949
rect 3603 1847 3637 1881
rect 3603 1779 3637 1813
rect 3603 1711 3637 1745
rect 3603 1643 3637 1677
rect 3603 1575 3637 1609
rect 3603 1507 3637 1541
rect 3603 1439 3637 1473
rect 3603 1371 3637 1405
rect 3603 1303 3637 1337
rect 3603 1235 3637 1269
rect 3603 1167 3637 1201
rect 3603 1099 3637 1133
rect 3603 1031 3637 1065
rect 3603 963 3637 997
rect 3603 895 3637 929
rect 3603 827 3637 861
rect 3603 759 3637 793
rect 3603 691 3637 725
rect 3603 623 3637 657
rect 3603 555 3637 589
rect 3603 487 3637 521
rect 3603 419 3637 453
rect 3603 351 3637 385
rect 3603 283 3637 317
rect 3603 215 3637 249
rect 3603 147 3637 181
rect 3603 79 3637 113
rect 3603 11 3637 45
rect 3603 -57 3637 -23
rect 3603 -125 3637 -91
rect 3603 -193 3637 -159
rect 3603 -261 3637 -227
rect 3603 -329 3637 -295
rect 3603 -397 3637 -363
rect 3603 -465 3637 -431
rect 3603 -533 3637 -499
rect -357 -567 -281 -533
rect -247 -567 -213 -533
rect -179 -567 -145 -533
rect -111 -567 -77 -533
rect -43 -567 -9 -533
rect 25 -567 59 -533
rect 93 -567 127 -533
rect 161 -567 195 -533
rect 229 -567 263 -533
rect 297 -567 331 -533
rect 365 -567 399 -533
rect 433 -567 467 -533
rect 501 -567 535 -533
rect 569 -567 603 -533
rect 637 -567 671 -533
rect 705 -567 739 -533
rect 773 -567 807 -533
rect 841 -567 875 -533
rect 909 -567 943 -533
rect 977 -567 1011 -533
rect 1045 -567 1079 -533
rect 1113 -567 1147 -533
rect 1181 -567 1215 -533
rect 1249 -567 1283 -533
rect 1317 -567 1351 -533
rect 1385 -567 1419 -533
rect 1453 -567 1487 -533
rect 1521 -567 1555 -533
rect 1589 -567 1623 -533
rect 1657 -567 1691 -533
rect 1725 -567 1759 -533
rect 1793 -567 1827 -533
rect 1861 -567 1895 -533
rect 1929 -567 1963 -533
rect 1997 -567 2031 -533
rect 2065 -567 2099 -533
rect 2133 -567 2167 -533
rect 2201 -567 2235 -533
rect 2269 -567 2303 -533
rect 2337 -567 2371 -533
rect 2405 -567 2439 -533
rect 2473 -567 2507 -533
rect 2541 -567 2575 -533
rect 2609 -567 2643 -533
rect 2677 -567 2711 -533
rect 2745 -567 2779 -533
rect 2813 -567 2847 -533
rect 2881 -567 2915 -533
rect 2949 -567 2983 -533
rect 3017 -567 3051 -533
rect 3085 -567 3119 -533
rect 3153 -567 3187 -533
rect 3221 -567 3255 -533
rect 3289 -567 3323 -533
rect 3357 -567 3391 -533
rect 3425 -567 3459 -533
rect 3493 -567 3527 -533
rect 3561 -567 3637 -533
<< metal1 >>
rect 3310 9486 3410 9510
rect 3310 9434 3334 9486
rect 3386 9434 3410 9486
rect 0 9200 3270 9260
rect 130 9100 3270 9200
rect 0 9040 3270 9100
rect 0 8840 190 9040
rect 360 8996 520 9010
rect 360 8944 374 8996
rect 426 8944 454 8996
rect 506 8944 520 8996
rect 360 8930 520 8944
rect 640 8996 800 9010
rect 640 8944 654 8996
rect 706 8944 734 8996
rect 786 8944 800 8996
rect 640 8930 800 8944
rect 920 8996 1080 9010
rect 920 8944 934 8996
rect 986 8944 1014 8996
rect 1066 8944 1080 8996
rect 920 8930 1080 8944
rect 1200 8996 1360 9010
rect 1200 8944 1214 8996
rect 1266 8944 1294 8996
rect 1346 8944 1360 8996
rect 1200 8930 1360 8944
rect 1480 8996 1640 9010
rect 1480 8944 1494 8996
rect 1546 8944 1574 8996
rect 1626 8944 1640 8996
rect 1480 8930 1640 8944
rect 1760 8996 1920 9010
rect 1760 8944 1774 8996
rect 1826 8944 1854 8996
rect 1906 8944 1920 8996
rect 1760 8930 1920 8944
rect 2040 8996 2200 9010
rect 2040 8944 2054 8996
rect 2106 8944 2134 8996
rect 2186 8944 2200 8996
rect 2040 8930 2200 8944
rect 2320 8996 2480 9010
rect 2320 8944 2334 8996
rect 2386 8944 2414 8996
rect 2466 8944 2480 8996
rect 2320 8930 2480 8944
rect 2600 8996 2760 9010
rect 2600 8944 2614 8996
rect 2666 8944 2694 8996
rect 2746 8944 2760 8996
rect 2600 8930 2760 8944
rect 2880 8996 3040 9010
rect 2880 8944 2894 8996
rect 2946 8944 2974 8996
rect 3026 8944 3040 8996
rect 2880 8930 3040 8944
rect 290 8896 380 8900
rect 290 8844 309 8896
rect 361 8844 380 8896
rect 290 8840 380 8844
rect 130 6840 190 8840
rect 410 7130 470 8930
rect 570 8896 660 8900
rect 570 8844 589 8896
rect 641 8844 660 8896
rect 570 8840 660 8844
rect 690 7130 750 8930
rect 850 8896 940 8900
rect 850 8844 869 8896
rect 921 8844 940 8896
rect 850 8840 940 8844
rect 970 7130 1030 8930
rect 1130 8896 1220 8900
rect 1130 8844 1149 8896
rect 1201 8844 1220 8896
rect 1130 8840 1220 8844
rect 1250 7130 1310 8930
rect 1410 8896 1500 8900
rect 1410 8844 1429 8896
rect 1481 8844 1500 8896
rect 1410 8840 1500 8844
rect 1530 7130 1590 8930
rect 1690 8896 1780 8900
rect 1690 8844 1709 8896
rect 1761 8844 1780 8896
rect 1690 8840 1780 8844
rect 1810 7130 1870 8930
rect 1970 8896 2060 8900
rect 1970 8844 1989 8896
rect 2041 8844 2060 8896
rect 1970 8840 2060 8844
rect 2090 7130 2150 8930
rect 2250 8896 2340 8900
rect 2250 8844 2269 8896
rect 2321 8844 2340 8896
rect 2250 8840 2340 8844
rect 2370 7130 2430 8930
rect 2530 8896 2620 8900
rect 2530 8844 2549 8896
rect 2601 8844 2620 8896
rect 2530 8840 2620 8844
rect 2650 7130 2710 8930
rect 2810 8896 2900 8900
rect 2810 8844 2829 8896
rect 2881 8844 2900 8896
rect 2810 8840 2900 8844
rect 2930 7130 2990 8930
rect 3080 8840 3270 9040
rect 3210 6840 3270 8840
rect 0 6580 190 6840
rect 290 6836 380 6840
rect 290 6784 309 6836
rect 361 6784 380 6836
rect 290 6780 380 6784
rect 570 6836 660 6840
rect 570 6784 589 6836
rect 641 6784 660 6836
rect 570 6780 660 6784
rect 850 6836 940 6840
rect 850 6784 869 6836
rect 921 6784 940 6836
rect 850 6780 940 6784
rect 1130 6836 1220 6840
rect 1130 6784 1149 6836
rect 1201 6784 1220 6836
rect 1130 6780 1220 6784
rect 1410 6836 1500 6840
rect 1410 6784 1429 6836
rect 1481 6784 1500 6836
rect 1410 6780 1500 6784
rect 1690 6836 1780 6840
rect 1690 6784 1709 6836
rect 1761 6784 1780 6836
rect 1690 6780 1780 6784
rect 1970 6836 2060 6840
rect 1970 6784 1989 6836
rect 2041 6784 2060 6836
rect 1970 6780 2060 6784
rect 2250 6836 2340 6840
rect 2250 6784 2269 6836
rect 2321 6784 2340 6836
rect 2250 6780 2340 6784
rect 2530 6836 2620 6840
rect 2530 6784 2549 6836
rect 2601 6784 2620 6836
rect 2530 6780 2620 6784
rect 2810 6836 2900 6840
rect 2810 6784 2829 6836
rect 2881 6784 2900 6836
rect 2810 6780 2900 6784
rect 360 6736 520 6750
rect 360 6684 374 6736
rect 426 6684 454 6736
rect 506 6684 520 6736
rect 360 6670 520 6684
rect 640 6736 800 6750
rect 640 6684 654 6736
rect 706 6684 734 6736
rect 786 6684 800 6736
rect 640 6670 800 6684
rect 920 6736 1080 6750
rect 920 6684 934 6736
rect 986 6684 1014 6736
rect 1066 6684 1080 6736
rect 920 6670 1080 6684
rect 1200 6736 1360 6750
rect 1200 6684 1214 6736
rect 1266 6684 1294 6736
rect 1346 6684 1360 6736
rect 1200 6670 1360 6684
rect 1430 6736 1590 6750
rect 1430 6684 1444 6736
rect 1496 6684 1524 6736
rect 1576 6684 1590 6736
rect 1430 6670 1590 6684
rect 290 6636 380 6640
rect 290 6584 309 6636
rect 361 6584 380 6636
rect 290 6580 380 6584
rect 130 4580 190 6580
rect 410 4870 470 6670
rect 570 6636 660 6640
rect 570 6584 589 6636
rect 641 6584 660 6636
rect 570 6580 660 6584
rect 690 4870 750 6670
rect 850 6636 940 6640
rect 850 6584 869 6636
rect 921 6584 940 6636
rect 850 6580 940 6584
rect 970 4870 1030 6670
rect 1130 6636 1220 6640
rect 1130 6584 1149 6636
rect 1201 6584 1220 6636
rect 1130 6580 1220 6584
rect 1250 4870 1310 6670
rect 1410 6636 1500 6640
rect 1410 6584 1429 6636
rect 1481 6584 1500 6636
rect 1410 6580 1500 6584
rect 1530 4950 1590 6670
rect 1810 6736 1970 6750
rect 1810 6684 1824 6736
rect 1876 6684 1904 6736
rect 1956 6684 1970 6736
rect 1810 6670 1970 6684
rect 2040 6736 2200 6750
rect 2040 6684 2054 6736
rect 2106 6684 2134 6736
rect 2186 6684 2200 6736
rect 2040 6670 2200 6684
rect 2320 6736 2480 6750
rect 2320 6684 2334 6736
rect 2386 6684 2414 6736
rect 2466 6684 2480 6736
rect 2320 6670 2480 6684
rect 2600 6736 2760 6750
rect 2600 6684 2614 6736
rect 2666 6684 2694 6736
rect 2746 6684 2760 6736
rect 2600 6670 2760 6684
rect 2830 6736 2990 6750
rect 2830 6684 2844 6736
rect 2896 6684 2924 6736
rect 2976 6684 2990 6736
rect 2830 6670 2990 6684
rect 1690 6636 1780 6640
rect 1690 6584 1709 6636
rect 1761 6584 1780 6636
rect 1690 6580 1780 6584
rect 1510 4936 1590 4950
rect 1510 4884 1524 4936
rect 1576 4884 1590 4936
rect 1510 4846 1590 4884
rect 1510 4794 1524 4846
rect 1576 4794 1590 4846
rect 1510 4780 1590 4794
rect 1810 4936 1870 6670
rect 1970 6636 2060 6640
rect 1970 6584 1989 6636
rect 2041 6584 2060 6636
rect 1970 6580 2060 6584
rect 1810 4884 1814 4936
rect 1866 4884 1870 4936
rect 1810 4856 1870 4884
rect 2090 4870 2150 6670
rect 2250 6636 2340 6640
rect 2250 6584 2269 6636
rect 2321 6584 2340 6636
rect 2250 6580 2340 6584
rect 2370 4870 2430 6670
rect 2530 6636 2620 6640
rect 2530 6584 2549 6636
rect 2601 6584 2620 6636
rect 2530 6580 2620 6584
rect 2650 4870 2710 6670
rect 2810 6636 2900 6640
rect 2810 6584 2829 6636
rect 2881 6584 2900 6636
rect 2810 6580 2900 6584
rect 2930 4870 2990 6670
rect 3080 6580 3270 6840
rect 1810 4804 1814 4856
rect 1866 4804 1870 4856
rect 1810 4790 1870 4804
rect 3210 4580 3270 6580
rect 0 4320 190 4580
rect 290 4576 380 4580
rect 290 4524 309 4576
rect 361 4524 380 4576
rect 290 4520 380 4524
rect 570 4576 660 4580
rect 570 4524 589 4576
rect 641 4524 660 4576
rect 570 4520 660 4524
rect 850 4576 940 4580
rect 850 4524 869 4576
rect 921 4524 940 4576
rect 850 4520 940 4524
rect 1130 4576 1220 4580
rect 1130 4524 1149 4576
rect 1201 4524 1220 4576
rect 1130 4520 1220 4524
rect 1410 4576 1500 4580
rect 1410 4524 1429 4576
rect 1481 4524 1500 4576
rect 1410 4520 1500 4524
rect 1690 4576 2060 4580
rect 1690 4524 1989 4576
rect 2041 4524 2060 4576
rect 1690 4520 2060 4524
rect 2250 4576 2340 4580
rect 2250 4524 2269 4576
rect 2321 4524 2340 4576
rect 2250 4520 2340 4524
rect 2530 4576 2620 4580
rect 2530 4524 2549 4576
rect 2601 4524 2620 4576
rect 2530 4520 2620 4524
rect 2810 4576 2900 4580
rect 2810 4524 2829 4576
rect 2881 4524 2900 4576
rect 2810 4520 2900 4524
rect 410 4476 570 4490
rect 410 4424 424 4476
rect 476 4424 504 4476
rect 556 4424 570 4476
rect 410 4410 570 4424
rect 640 4476 800 4490
rect 640 4424 654 4476
rect 706 4424 734 4476
rect 786 4424 800 4476
rect 640 4410 800 4424
rect 920 4476 1080 4490
rect 920 4424 934 4476
rect 986 4424 1014 4476
rect 1066 4424 1080 4476
rect 920 4410 1080 4424
rect 1200 4476 1360 4490
rect 1200 4424 1214 4476
rect 1266 4424 1294 4476
rect 1346 4424 1360 4476
rect 1200 4410 1360 4424
rect 1430 4476 1590 4490
rect 1430 4424 1444 4476
rect 1496 4424 1524 4476
rect 1576 4424 1590 4476
rect 1430 4410 1590 4424
rect 290 4376 380 4380
rect 290 4324 309 4376
rect 361 4324 380 4376
rect 290 4320 380 4324
rect 130 2320 190 4320
rect 410 2610 470 4410
rect 570 4376 660 4380
rect 570 4324 589 4376
rect 641 4324 660 4376
rect 570 4320 660 4324
rect 690 2610 750 4410
rect 850 4376 940 4380
rect 850 4324 869 4376
rect 921 4324 940 4376
rect 850 4320 940 4324
rect 970 2610 1030 4410
rect 1130 4376 1220 4380
rect 1130 4324 1149 4376
rect 1201 4324 1220 4376
rect 1130 4320 1220 4324
rect 1250 2610 1310 4410
rect 1410 4376 1500 4380
rect 1410 4324 1429 4376
rect 1481 4324 1500 4376
rect 1410 4320 1500 4324
rect 1530 2610 1590 4410
rect 1810 4476 2200 4490
rect 1810 4424 2049 4476
rect 2101 4424 2134 4476
rect 2186 4424 2200 4476
rect 1810 4410 2200 4424
rect 2320 4476 2480 4490
rect 2320 4424 2334 4476
rect 2386 4424 2414 4476
rect 2466 4424 2480 4476
rect 2320 4410 2480 4424
rect 2600 4476 2760 4490
rect 2600 4424 2614 4476
rect 2666 4424 2694 4476
rect 2746 4424 2760 4476
rect 2600 4410 2760 4424
rect 2830 4476 2990 4490
rect 2830 4424 2844 4476
rect 2896 4424 2924 4476
rect 2976 4424 2990 4476
rect 2830 4410 2990 4424
rect 1690 4376 1780 4380
rect 1690 4324 1709 4376
rect 1761 4324 1780 4376
rect 1690 4320 1780 4324
rect 1810 2610 1870 4410
rect 1970 4376 2060 4380
rect 1970 4324 1989 4376
rect 2041 4324 2060 4376
rect 1970 4320 2060 4324
rect 2090 2610 2150 4410
rect 2250 4376 2340 4380
rect 2250 4324 2269 4376
rect 2321 4324 2340 4376
rect 2250 4320 2340 4324
rect 2370 2610 2430 4410
rect 2530 4376 2620 4380
rect 2530 4324 2549 4376
rect 2601 4324 2620 4376
rect 2530 4320 2620 4324
rect 2650 2610 2710 4410
rect 2810 4376 2900 4380
rect 2810 4324 2829 4376
rect 2881 4324 2900 4376
rect 2810 4320 2900 4324
rect 2930 2610 2990 4410
rect 3080 4320 3270 4580
rect 3310 6726 3410 9434
rect 3310 6674 3334 6726
rect 3386 6674 3410 6726
rect 3310 6646 3410 6674
rect 3310 6594 3334 6646
rect 3386 6594 3410 6646
rect 3310 4466 3410 6594
rect 3310 4414 3334 4466
rect 3386 4414 3410 4466
rect 3310 4386 3410 4414
rect 3310 4334 3334 4386
rect 3386 4334 3410 4386
rect 3310 4320 3410 4334
rect 3210 2320 3270 4320
rect 0 2060 190 2320
rect 290 2316 380 2320
rect 290 2264 309 2316
rect 361 2264 380 2316
rect 290 2260 380 2264
rect 570 2316 660 2320
rect 570 2264 589 2316
rect 641 2264 660 2316
rect 570 2260 660 2264
rect 850 2316 940 2320
rect 850 2264 869 2316
rect 921 2264 940 2316
rect 850 2260 940 2264
rect 1130 2316 1220 2320
rect 1130 2264 1149 2316
rect 1201 2264 1220 2316
rect 1130 2260 1220 2264
rect 1410 2316 1500 2320
rect 1410 2264 1429 2316
rect 1481 2264 1500 2316
rect 1410 2260 1500 2264
rect 1690 2316 1780 2320
rect 1690 2264 1709 2316
rect 1761 2264 1780 2316
rect 1690 2260 1780 2264
rect 1970 2316 2060 2320
rect 1970 2264 1989 2316
rect 2041 2264 2060 2316
rect 1970 2260 2060 2264
rect 2250 2316 2340 2320
rect 2250 2264 2269 2316
rect 2321 2264 2340 2316
rect 2250 2260 2340 2264
rect 2530 2316 2620 2320
rect 2530 2264 2549 2316
rect 2601 2264 2620 2316
rect 2530 2260 2620 2264
rect 2810 2316 2900 2320
rect 2810 2264 2829 2316
rect 2881 2264 2900 2316
rect 2810 2260 2900 2264
rect 410 2216 570 2230
rect 410 2164 424 2216
rect 476 2164 504 2216
rect 556 2164 570 2216
rect 410 2150 570 2164
rect 640 2216 800 2230
rect 640 2164 654 2216
rect 706 2164 734 2216
rect 786 2164 800 2216
rect 640 2150 800 2164
rect 920 2216 1080 2230
rect 920 2164 934 2216
rect 986 2164 1014 2216
rect 1066 2164 1080 2216
rect 920 2150 1080 2164
rect 1200 2216 1360 2230
rect 1200 2164 1214 2216
rect 1266 2164 1294 2216
rect 1346 2164 1360 2216
rect 1200 2150 1360 2164
rect 1430 2216 1590 2230
rect 1430 2164 1444 2216
rect 1496 2164 1524 2216
rect 1576 2164 1590 2216
rect 1430 2150 1590 2164
rect 290 2116 380 2120
rect 290 2064 309 2116
rect 361 2064 380 2116
rect 290 2060 380 2064
rect 130 60 190 2060
rect 410 350 470 2150
rect 570 2116 660 2120
rect 570 2064 589 2116
rect 641 2064 660 2116
rect 570 2060 660 2064
rect 690 350 750 2150
rect 850 2116 940 2120
rect 850 2064 869 2116
rect 921 2064 940 2116
rect 850 2060 940 2064
rect 970 350 1030 2150
rect 1130 2116 1220 2120
rect 1130 2064 1149 2116
rect 1201 2064 1220 2116
rect 1130 2060 1220 2064
rect 1250 350 1310 2150
rect 1410 2116 1500 2120
rect 1410 2064 1429 2116
rect 1481 2064 1500 2116
rect 1410 2060 1500 2064
rect 1530 350 1590 2150
rect 1810 2216 1970 2230
rect 1810 2164 1824 2216
rect 1876 2164 1904 2216
rect 1956 2164 1970 2216
rect 1810 2150 1970 2164
rect 2040 2216 2200 2230
rect 2040 2164 2054 2216
rect 2106 2164 2134 2216
rect 2186 2164 2200 2216
rect 2040 2150 2200 2164
rect 2320 2216 2480 2230
rect 2320 2164 2334 2216
rect 2386 2164 2414 2216
rect 2466 2164 2480 2216
rect 2320 2150 2480 2164
rect 2600 2216 2760 2230
rect 2600 2164 2614 2216
rect 2666 2164 2694 2216
rect 2746 2164 2760 2216
rect 2600 2150 2760 2164
rect 2830 2216 2990 2230
rect 2830 2164 2844 2216
rect 2896 2164 2924 2216
rect 2976 2164 2990 2216
rect 2830 2150 2990 2164
rect 1690 2116 1780 2120
rect 1690 2064 1709 2116
rect 1761 2064 1780 2116
rect 1690 2060 1780 2064
rect 1810 350 1870 2150
rect 1970 2116 2060 2120
rect 1970 2064 1989 2116
rect 2041 2064 2060 2116
rect 1970 2060 2060 2064
rect 2090 350 2150 2150
rect 2250 2116 2340 2120
rect 2250 2064 2269 2116
rect 2321 2064 2340 2116
rect 2250 2060 2340 2064
rect 2370 350 2430 2150
rect 2530 2116 2620 2120
rect 2530 2064 2549 2116
rect 2601 2064 2620 2116
rect 2530 2060 2620 2064
rect 2650 350 2710 2150
rect 2810 2116 2900 2120
rect 2810 2064 2829 2116
rect 2881 2064 2900 2116
rect 2810 2060 2900 2064
rect 2930 350 2990 2150
rect 3070 2060 3270 2320
rect 3210 60 3270 2060
rect 0 -60 190 60
rect 290 56 380 60
rect 290 4 309 56
rect 361 4 380 56
rect 290 0 380 4
rect 570 56 660 60
rect 570 4 589 56
rect 641 4 660 56
rect 570 0 660 4
rect 850 56 940 60
rect 850 4 869 56
rect 921 4 940 56
rect 850 0 940 4
rect 1130 56 1220 60
rect 1130 4 1149 56
rect 1201 4 1220 56
rect 1130 0 1220 4
rect 1410 56 1500 60
rect 1410 4 1429 56
rect 1481 4 1500 56
rect 1410 0 1500 4
rect 1690 56 1780 60
rect 1690 4 1709 56
rect 1761 4 1780 56
rect 1690 0 1780 4
rect 1970 56 2060 60
rect 1970 4 1989 56
rect 2041 4 2060 56
rect 1970 0 2060 4
rect 2250 56 2340 60
rect 2250 4 2269 56
rect 2321 4 2340 56
rect 2250 0 2340 4
rect 2530 56 2620 60
rect 2530 4 2549 56
rect 2601 4 2620 56
rect 2530 0 2620 4
rect 2810 56 2900 60
rect 2810 4 2829 56
rect 2881 4 2900 56
rect 2810 0 2900 4
rect 3080 -60 3270 60
rect 0 -120 3270 -60
rect 130 -220 3270 -120
rect 0 -280 3270 -220
rect 3310 2396 3390 2400
rect 3310 2344 3324 2396
rect 3376 2344 3390 2396
rect 3310 2316 3390 2344
rect 3310 2264 3324 2316
rect 3376 2264 3390 2316
rect 3310 136 3390 2264
rect 3310 84 3324 136
rect 3376 84 3390 136
rect 3310 56 3390 84
rect 3310 4 3324 56
rect 3376 4 3390 56
rect 3310 -310 3390 4
rect 3220 -324 3390 -310
rect 3220 -376 3234 -324
rect 3286 -376 3324 -324
rect 3376 -376 3390 -324
rect 3220 -390 3390 -376
<< via1 >>
rect 3334 9434 3386 9486
rect 374 8944 426 8996
rect 454 8944 506 8996
rect 654 8944 706 8996
rect 734 8944 786 8996
rect 934 8944 986 8996
rect 1014 8944 1066 8996
rect 1214 8944 1266 8996
rect 1294 8944 1346 8996
rect 1494 8944 1546 8996
rect 1574 8944 1626 8996
rect 1774 8944 1826 8996
rect 1854 8944 1906 8996
rect 2054 8944 2106 8996
rect 2134 8944 2186 8996
rect 2334 8944 2386 8996
rect 2414 8944 2466 8996
rect 2614 8944 2666 8996
rect 2694 8944 2746 8996
rect 2894 8944 2946 8996
rect 2974 8944 3026 8996
rect 309 8844 361 8896
rect 589 8844 641 8896
rect 869 8844 921 8896
rect 1149 8844 1201 8896
rect 1429 8844 1481 8896
rect 1709 8844 1761 8896
rect 1989 8844 2041 8896
rect 2269 8844 2321 8896
rect 2549 8844 2601 8896
rect 2829 8844 2881 8896
rect 309 6784 361 6836
rect 589 6784 641 6836
rect 869 6784 921 6836
rect 1149 6784 1201 6836
rect 1429 6784 1481 6836
rect 1709 6784 1761 6836
rect 1989 6784 2041 6836
rect 2269 6784 2321 6836
rect 2549 6784 2601 6836
rect 2829 6784 2881 6836
rect 374 6684 426 6736
rect 454 6684 506 6736
rect 654 6684 706 6736
rect 734 6684 786 6736
rect 934 6684 986 6736
rect 1014 6684 1066 6736
rect 1214 6684 1266 6736
rect 1294 6684 1346 6736
rect 1444 6684 1496 6736
rect 1524 6684 1576 6736
rect 309 6584 361 6636
rect 589 6584 641 6636
rect 869 6584 921 6636
rect 1149 6584 1201 6636
rect 1429 6584 1481 6636
rect 1824 6684 1876 6736
rect 1904 6684 1956 6736
rect 2054 6684 2106 6736
rect 2134 6684 2186 6736
rect 2334 6684 2386 6736
rect 2414 6684 2466 6736
rect 2614 6684 2666 6736
rect 2694 6684 2746 6736
rect 2844 6684 2896 6736
rect 2924 6684 2976 6736
rect 1709 6584 1761 6636
rect 1524 4884 1576 4936
rect 1524 4794 1576 4846
rect 1989 6584 2041 6636
rect 1814 4884 1866 4936
rect 2269 6584 2321 6636
rect 2549 6584 2601 6636
rect 2829 6584 2881 6636
rect 1814 4804 1866 4856
rect 309 4524 361 4576
rect 589 4524 641 4576
rect 869 4524 921 4576
rect 1149 4524 1201 4576
rect 1429 4524 1481 4576
rect 1989 4524 2041 4576
rect 2269 4524 2321 4576
rect 2549 4524 2601 4576
rect 2829 4524 2881 4576
rect 424 4424 476 4476
rect 504 4424 556 4476
rect 654 4424 706 4476
rect 734 4424 786 4476
rect 934 4424 986 4476
rect 1014 4424 1066 4476
rect 1214 4424 1266 4476
rect 1294 4424 1346 4476
rect 1444 4424 1496 4476
rect 1524 4424 1576 4476
rect 309 4324 361 4376
rect 589 4324 641 4376
rect 869 4324 921 4376
rect 1149 4324 1201 4376
rect 1429 4324 1481 4376
rect 2049 4424 2101 4476
rect 2134 4424 2186 4476
rect 2334 4424 2386 4476
rect 2414 4424 2466 4476
rect 2614 4424 2666 4476
rect 2694 4424 2746 4476
rect 2844 4424 2896 4476
rect 2924 4424 2976 4476
rect 1709 4324 1761 4376
rect 1989 4324 2041 4376
rect 2269 4324 2321 4376
rect 2549 4324 2601 4376
rect 2829 4324 2881 4376
rect 3334 6674 3386 6726
rect 3334 6594 3386 6646
rect 3334 4414 3386 4466
rect 3334 4334 3386 4386
rect 309 2264 361 2316
rect 589 2264 641 2316
rect 869 2264 921 2316
rect 1149 2264 1201 2316
rect 1429 2264 1481 2316
rect 1709 2264 1761 2316
rect 1989 2264 2041 2316
rect 2269 2264 2321 2316
rect 2549 2264 2601 2316
rect 2829 2264 2881 2316
rect 424 2164 476 2216
rect 504 2164 556 2216
rect 654 2164 706 2216
rect 734 2164 786 2216
rect 934 2164 986 2216
rect 1014 2164 1066 2216
rect 1214 2164 1266 2216
rect 1294 2164 1346 2216
rect 1444 2164 1496 2216
rect 1524 2164 1576 2216
rect 309 2064 361 2116
rect 589 2064 641 2116
rect 869 2064 921 2116
rect 1149 2064 1201 2116
rect 1429 2064 1481 2116
rect 1824 2164 1876 2216
rect 1904 2164 1956 2216
rect 2054 2164 2106 2216
rect 2134 2164 2186 2216
rect 2334 2164 2386 2216
rect 2414 2164 2466 2216
rect 2614 2164 2666 2216
rect 2694 2164 2746 2216
rect 2844 2164 2896 2216
rect 2924 2164 2976 2216
rect 1709 2064 1761 2116
rect 1989 2064 2041 2116
rect 2269 2064 2321 2116
rect 2549 2064 2601 2116
rect 2829 2064 2881 2116
rect 309 4 361 56
rect 589 4 641 56
rect 869 4 921 56
rect 1149 4 1201 56
rect 1429 4 1481 56
rect 1709 4 1761 56
rect 1989 4 2041 56
rect 2269 4 2321 56
rect 2549 4 2601 56
rect 2829 4 2881 56
rect 3324 2344 3376 2396
rect 3324 2264 3376 2316
rect 3324 84 3376 136
rect 3324 4 3376 56
rect 3234 -376 3286 -324
rect 3324 -376 3376 -324
<< metal2 >>
rect 3310 9488 3410 9510
rect 3310 9432 3332 9488
rect 3388 9432 3410 9488
rect 3310 9410 3410 9432
rect 360 8998 3410 9010
rect 360 8996 3237 8998
rect 360 8944 374 8996
rect 426 8944 454 8996
rect 506 8944 654 8996
rect 706 8944 734 8996
rect 786 8944 934 8996
rect 986 8944 1014 8996
rect 1066 8944 1214 8996
rect 1266 8944 1294 8996
rect 1346 8944 1494 8996
rect 1546 8944 1574 8996
rect 1626 8944 1774 8996
rect 1826 8944 1854 8996
rect 1906 8944 2054 8996
rect 2106 8944 2134 8996
rect 2186 8944 2334 8996
rect 2386 8944 2414 8996
rect 2466 8944 2614 8996
rect 2666 8944 2694 8996
rect 2746 8944 2894 8996
rect 2946 8944 2974 8996
rect 3026 8944 3237 8996
rect 360 8942 3237 8944
rect 3293 8942 3337 8998
rect 3393 8942 3410 8998
rect 360 8930 3410 8942
rect -130 8896 3470 8900
rect -130 8888 309 8896
rect -130 8832 -108 8888
rect -52 8844 309 8888
rect 361 8844 589 8896
rect 641 8844 869 8896
rect 921 8844 1149 8896
rect 1201 8844 1429 8896
rect 1481 8844 1709 8896
rect 1761 8844 1989 8896
rect 2041 8844 2269 8896
rect 2321 8844 2549 8896
rect 2601 8844 2829 8896
rect 2881 8844 3470 8896
rect -52 8840 3470 8844
rect -52 8832 -30 8840
rect -130 8798 -30 8832
rect -130 8742 -108 8798
rect -52 8742 -30 8798
rect -130 8730 -30 8742
rect -290 6938 -190 6950
rect -290 6882 -268 6938
rect -212 6882 -190 6938
rect -290 6848 -190 6882
rect -290 6792 -268 6848
rect -212 6840 -190 6848
rect -212 6836 1510 6840
rect -212 6792 309 6836
rect -290 6784 309 6792
rect 361 6784 589 6836
rect 641 6784 869 6836
rect 921 6784 1149 6836
rect 1201 6784 1429 6836
rect 1481 6784 1510 6836
rect -290 6780 1510 6784
rect 1690 6836 3570 6840
rect 1690 6784 1709 6836
rect 1761 6784 1989 6836
rect 2041 6784 2269 6836
rect 2321 6784 2549 6836
rect 2601 6784 2829 6836
rect 2881 6828 3570 6836
rect 2881 6784 3492 6828
rect 1690 6780 3492 6784
rect 3470 6772 3492 6780
rect 3548 6772 3570 6828
rect -510 6750 -410 6760
rect -510 6738 1590 6750
rect -510 6682 -488 6738
rect -432 6736 1590 6738
rect -432 6684 374 6736
rect 426 6684 454 6736
rect 506 6684 654 6736
rect 706 6684 734 6736
rect 786 6684 934 6736
rect 986 6684 1014 6736
rect 1066 6684 1214 6736
rect 1266 6684 1294 6736
rect 1346 6684 1444 6736
rect 1496 6684 1524 6736
rect 1576 6684 1590 6736
rect -432 6682 1590 6684
rect -510 6670 1590 6682
rect 1810 6736 2990 6750
rect 1810 6684 1824 6736
rect 1876 6684 1904 6736
rect 1956 6684 2054 6736
rect 2106 6684 2134 6736
rect 2186 6684 2334 6736
rect 2386 6684 2414 6736
rect 2466 6684 2614 6736
rect 2666 6684 2694 6736
rect 2746 6684 2844 6736
rect 2896 6684 2924 6736
rect 2976 6684 2990 6736
rect 1810 6670 2990 6684
rect 3310 6726 3410 6740
rect 3310 6674 3334 6726
rect 3386 6674 3410 6726
rect -510 6660 -410 6670
rect 3310 6646 3410 6674
rect 3470 6738 3570 6772
rect 3470 6682 3492 6738
rect 3548 6682 3570 6738
rect 3470 6670 3570 6682
rect 3310 6640 3334 6646
rect 290 6636 3334 6640
rect 290 6584 309 6636
rect 361 6584 589 6636
rect 641 6584 869 6636
rect 921 6584 1149 6636
rect 1201 6584 1429 6636
rect 1481 6584 1709 6636
rect 1761 6584 1989 6636
rect 2041 6584 2269 6636
rect 2321 6584 2549 6636
rect 2601 6584 2829 6636
rect 2881 6594 3334 6636
rect 3386 6594 3410 6646
rect 2881 6584 3410 6594
rect 290 6580 3410 6584
rect 1510 4938 1590 4950
rect 1510 4882 1522 4938
rect 1578 4882 1590 4938
rect 1510 4848 1590 4882
rect 1510 4792 1522 4848
rect 1578 4792 1590 4848
rect 1510 4780 1590 4792
rect 1810 4936 1870 4950
rect 1810 4884 1814 4936
rect 1866 4884 1870 4936
rect 1810 4856 1870 4884
rect 1810 4804 1814 4856
rect 1866 4804 1870 4856
rect -290 4678 -190 4690
rect -290 4622 -268 4678
rect -212 4622 -190 4678
rect -290 4588 -190 4622
rect -290 4532 -268 4588
rect -212 4580 -190 4588
rect -212 4576 1510 4580
rect -212 4532 309 4576
rect -290 4524 309 4532
rect 361 4524 589 4576
rect 641 4524 869 4576
rect 921 4524 1149 4576
rect 1201 4524 1429 4576
rect 1481 4524 1510 4576
rect -290 4520 1510 4524
rect -510 4490 -410 4500
rect 1810 4490 1870 4804
rect 3470 4678 3570 4690
rect 3470 4622 3492 4678
rect 3548 4622 3570 4678
rect 3470 4588 3570 4622
rect 3470 4580 3492 4588
rect 1970 4576 3492 4580
rect 1970 4524 1989 4576
rect 2041 4524 2269 4576
rect 2321 4524 2549 4576
rect 2601 4524 2829 4576
rect 2881 4532 3492 4576
rect 3548 4532 3570 4588
rect 2881 4524 3570 4532
rect 1970 4520 3570 4524
rect -510 4478 1870 4490
rect -510 4422 -488 4478
rect -432 4476 1870 4478
rect -432 4424 424 4476
rect 476 4424 504 4476
rect 556 4424 654 4476
rect 706 4424 734 4476
rect 786 4424 934 4476
rect 986 4424 1014 4476
rect 1066 4424 1214 4476
rect 1266 4424 1294 4476
rect 1346 4424 1444 4476
rect 1496 4424 1524 4476
rect 1576 4424 1870 4476
rect -432 4422 1870 4424
rect -510 4410 1870 4422
rect 2040 4478 2990 4490
rect 2040 4422 2042 4478
rect 2098 4476 2132 4478
rect 2188 4476 2990 4478
rect 2101 4424 2132 4476
rect 2188 4424 2334 4476
rect 2386 4424 2414 4476
rect 2466 4424 2614 4476
rect 2666 4424 2694 4476
rect 2746 4424 2844 4476
rect 2896 4424 2924 4476
rect 2976 4424 2990 4476
rect 2098 4422 2132 4424
rect 2188 4422 2990 4424
rect 2040 4410 2990 4422
rect 3310 4466 3410 4480
rect 3310 4414 3334 4466
rect 3386 4414 3410 4466
rect -510 4400 -410 4410
rect 3310 4386 3410 4414
rect 3310 4380 3334 4386
rect 290 4376 3334 4380
rect 290 4324 309 4376
rect 361 4324 589 4376
rect 641 4324 869 4376
rect 921 4324 1149 4376
rect 1201 4324 1429 4376
rect 1481 4324 1709 4376
rect 1761 4324 1989 4376
rect 2041 4324 2269 4376
rect 2321 4324 2549 4376
rect 2601 4324 2829 4376
rect 2881 4334 3334 4376
rect 3386 4334 3410 4386
rect 2881 4324 3410 4334
rect 290 4320 3410 4324
rect 3310 2396 3390 2400
rect 3310 2344 3324 2396
rect 3376 2344 3390 2396
rect 3310 2320 3390 2344
rect -110 2316 1510 2320
rect -110 2264 309 2316
rect 361 2264 589 2316
rect 641 2264 869 2316
rect 921 2264 1149 2316
rect 1201 2264 1429 2316
rect 1481 2264 1510 2316
rect -110 2260 1510 2264
rect 1690 2316 3390 2320
rect 1690 2264 1709 2316
rect 1761 2264 1989 2316
rect 2041 2264 2269 2316
rect 2321 2264 2549 2316
rect 2601 2264 2829 2316
rect 2881 2264 3324 2316
rect 3376 2264 3390 2316
rect 1690 2260 3390 2264
rect -110 60 -30 2260
rect 3690 2230 3790 2240
rect 410 2218 3790 2230
rect 410 2216 3237 2218
rect 410 2164 424 2216
rect 476 2164 504 2216
rect 556 2164 654 2216
rect 706 2164 734 2216
rect 786 2164 934 2216
rect 986 2164 1014 2216
rect 1066 2164 1214 2216
rect 1266 2164 1294 2216
rect 1346 2164 1444 2216
rect 1496 2164 1524 2216
rect 1576 2164 1824 2216
rect 1876 2164 1904 2216
rect 1956 2164 2054 2216
rect 2106 2164 2134 2216
rect 2186 2164 2334 2216
rect 2386 2164 2414 2216
rect 2466 2164 2614 2216
rect 2666 2164 2694 2216
rect 2746 2164 2844 2216
rect 2896 2164 2924 2216
rect 2976 2164 3237 2216
rect 410 2162 3237 2164
rect 3293 2162 3337 2218
rect 3393 2162 3712 2218
rect 3768 2162 3790 2218
rect 410 2150 3790 2162
rect 3690 2140 3790 2150
rect 10 2128 300 2140
rect 10 2072 22 2128
rect 78 2072 112 2128
rect 168 2072 202 2128
rect 258 2120 300 2128
rect 258 2116 2910 2120
rect 258 2072 309 2116
rect 10 2064 309 2072
rect 361 2064 589 2116
rect 641 2064 869 2116
rect 921 2064 1149 2116
rect 1201 2064 1429 2116
rect 1481 2064 1709 2116
rect 1761 2064 1989 2116
rect 2041 2064 2269 2116
rect 2321 2064 2549 2116
rect 2601 2064 2829 2116
rect 2881 2064 2910 2116
rect 10 2060 2910 2064
rect 3310 136 3390 140
rect 3310 84 3324 136
rect 3376 84 3390 136
rect 3310 60 3390 84
rect -110 56 1500 60
rect -110 4 309 56
rect 361 4 589 56
rect 641 4 869 56
rect 921 4 1149 56
rect 1201 4 1429 56
rect 1481 4 1500 56
rect -110 0 1500 4
rect 1690 56 3390 60
rect 1690 4 1709 56
rect 1761 4 1989 56
rect 2041 4 2269 56
rect 2321 4 2549 56
rect 2601 4 2829 56
rect 2881 4 3324 56
rect 3376 4 3390 56
rect 1690 0 3390 4
rect -110 -420 -30 0
rect 20 -322 3390 -310
rect 20 -378 32 -322
rect 88 -378 122 -322
rect 178 -324 3390 -322
rect 178 -376 3234 -324
rect 3286 -376 3324 -324
rect 3376 -376 3390 -324
rect 178 -378 3390 -376
rect 20 -390 3390 -378
rect -110 -432 3570 -420
rect -110 -488 3392 -432
rect 3448 -488 3492 -432
rect 3548 -488 3570 -432
rect -110 -500 3570 -488
rect 20 -590 100 -500
rect 10 -612 110 -590
rect 10 -668 32 -612
rect 88 -668 110 -612
rect 10 -690 110 -668
<< via2 >>
rect 3332 9486 3388 9488
rect 3332 9434 3334 9486
rect 3334 9434 3386 9486
rect 3386 9434 3388 9486
rect 3332 9432 3388 9434
rect 3237 8942 3293 8998
rect 3337 8942 3393 8998
rect -108 8832 -52 8888
rect -108 8742 -52 8798
rect -268 6882 -212 6938
rect -268 6792 -212 6848
rect 3492 6772 3548 6828
rect -488 6682 -432 6738
rect 3492 6682 3548 6738
rect 1522 4936 1578 4938
rect 1522 4884 1524 4936
rect 1524 4884 1576 4936
rect 1576 4884 1578 4936
rect 1522 4882 1578 4884
rect 1522 4846 1578 4848
rect 1522 4794 1524 4846
rect 1524 4794 1576 4846
rect 1576 4794 1578 4846
rect 1522 4792 1578 4794
rect -268 4622 -212 4678
rect -268 4532 -212 4588
rect 3492 4622 3548 4678
rect 3492 4532 3548 4588
rect -488 4422 -432 4478
rect 2042 4476 2098 4478
rect 2132 4476 2188 4478
rect 2042 4424 2049 4476
rect 2049 4424 2098 4476
rect 2132 4424 2134 4476
rect 2134 4424 2186 4476
rect 2186 4424 2188 4476
rect 2042 4422 2098 4424
rect 2132 4422 2188 4424
rect 3237 2162 3293 2218
rect 3337 2162 3393 2218
rect 3712 2162 3768 2218
rect 22 2072 78 2128
rect 112 2072 168 2128
rect 202 2072 258 2128
rect 32 -378 88 -322
rect 122 -378 178 -322
rect 3392 -488 3448 -432
rect 3492 -488 3548 -432
rect 32 -668 88 -612
<< metal3 >>
rect -130 8888 -30 9510
rect 3310 9488 3410 9510
rect 3310 9432 3332 9488
rect 3388 9432 3410 9488
rect 3310 9410 3410 9432
rect 3220 8998 3410 9010
rect 3220 8942 3237 8998
rect 3293 8942 3337 8998
rect 3393 8942 3410 8998
rect 3220 8930 3410 8942
rect -130 8832 -108 8888
rect -52 8832 -30 8888
rect -130 8798 -30 8832
rect -130 8742 -108 8798
rect -52 8742 -30 8798
rect -290 6938 -190 6950
rect -290 6882 -268 6938
rect -212 6882 -190 6938
rect -290 6848 -190 6882
rect -290 6792 -268 6848
rect -212 6792 -190 6848
rect -500 6738 -420 6750
rect -500 6682 -488 6738
rect -432 6682 -420 6738
rect -500 6670 -420 6682
rect -290 4678 -190 6792
rect -290 4622 -268 4678
rect -212 4622 -190 4678
rect -290 4588 -190 4622
rect -290 4532 -268 4588
rect -212 4532 -190 4588
rect -500 4478 -420 4490
rect -500 4422 -488 4478
rect -432 4422 -420 4478
rect -500 4410 -420 4422
rect -290 -310 -190 4532
rect -130 2140 -30 8742
rect 1510 4938 1590 4950
rect 1510 4882 1522 4938
rect 1578 4882 1590 4938
rect 1510 4848 1590 4882
rect 1510 4792 1522 4848
rect 1578 4792 1590 4848
rect 1510 4780 1590 4792
rect 1530 4490 1590 4780
rect 1530 4478 2200 4490
rect 1530 4422 2042 4478
rect 2098 4422 2132 4478
rect 2188 4422 2200 4478
rect 1530 4410 2200 4422
rect 3310 2230 3410 8930
rect 3220 2218 3410 2230
rect 3220 2162 3237 2218
rect 3293 2162 3337 2218
rect 3393 2162 3410 2218
rect 3220 2150 3410 2162
rect 3470 6828 3570 6840
rect 3470 6772 3492 6828
rect 3548 6772 3570 6828
rect 3470 6738 3570 6772
rect 3470 6682 3492 6738
rect 3548 6682 3570 6738
rect 3470 4678 3570 6682
rect 3470 4622 3492 4678
rect 3548 4622 3570 4678
rect 3470 4588 3570 4622
rect 3470 4532 3492 4588
rect 3548 4532 3570 4588
rect -130 2128 300 2140
rect -130 2072 22 2128
rect 78 2072 112 2128
rect 168 2072 202 2128
rect 258 2072 300 2128
rect -130 2060 300 2072
rect -290 -322 200 -310
rect -290 -378 32 -322
rect 88 -378 122 -322
rect 178 -378 200 -322
rect -290 -390 200 -378
rect -290 -690 -190 -390
rect 3470 -420 3570 4532
rect 3690 2218 3790 2240
rect 3690 2162 3712 2218
rect 3768 2162 3790 2218
rect 3690 2140 3790 2162
rect 3380 -432 3570 -420
rect 3380 -488 3392 -432
rect 3448 -488 3492 -432
rect 3548 -488 3570 -432
rect 3380 -500 3570 -488
rect 10 -612 110 -590
rect 10 -668 32 -612
rect 88 -668 110 -612
rect 10 -690 110 -668
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_0
timestamp 1757161594
transform 0 1 3167 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_1
timestamp 1757161594
transform 0 1 2607 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_2
timestamp 1757161594
transform 0 1 2887 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_3
timestamp 1757161594
transform 0 1 2327 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_4
timestamp 1757161594
transform 0 1 2047 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_5
timestamp 1757161594
transform 0 1 1767 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_6
timestamp 1757161594
transform 0 1 927 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_7
timestamp 1757161594
transform 0 1 1207 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_8
timestamp 1757161594
transform 0 1 1487 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_9
timestamp 1757161594
transform 0 1 647 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_10
timestamp 1757161594
transform 0 1 367 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_11
timestamp 1757161594
transform 0 1 87 1 0 1058
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_12
timestamp 1757161594
transform 0 1 3167 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_13
timestamp 1757161594
transform 0 1 2887 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_14
timestamp 1757161594
transform 0 1 2607 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_15
timestamp 1757161594
transform 0 1 2327 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_16
timestamp 1757161594
transform 0 1 2047 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_17
timestamp 1757161594
transform 0 1 1767 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_18
timestamp 1757161594
transform 0 1 1487 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_19
timestamp 1757161594
transform 0 1 1207 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_20
timestamp 1757161594
transform 0 1 927 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_21
timestamp 1757161594
transform 0 1 647 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_22
timestamp 1757161594
transform 0 1 367 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_23
timestamp 1757161594
transform 0 1 87 1 0 3318
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_24
timestamp 1757161594
transform 0 1 2887 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_25
timestamp 1757161594
transform 0 1 3167 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_26
timestamp 1757161594
transform 0 1 2327 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_27
timestamp 1757161594
transform 0 1 2607 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_28
timestamp 1757161594
transform 0 1 1767 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_29
timestamp 1757161594
transform 0 1 2047 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_30
timestamp 1757161594
transform 0 1 1207 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_31
timestamp 1757161594
transform 0 1 1487 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_32
timestamp 1757161594
transform 0 1 647 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_33
timestamp 1757161594
transform 0 1 927 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_34
timestamp 1757161594
transform 0 1 87 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_35
timestamp 1757161594
transform 0 1 367 1 0 5578
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_36
timestamp 1757161594
transform 0 1 647 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_37
timestamp 1757161594
transform 0 1 927 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_38
timestamp 1757161594
transform 0 1 87 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_39
timestamp 1757161594
transform 0 1 367 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_40
timestamp 1757161594
transform 0 1 2327 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_41
timestamp 1757161594
transform 0 1 1767 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_42
timestamp 1757161594
transform 0 1 2047 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_43
timestamp 1757161594
transform 0 1 1207 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_44
timestamp 1757161594
transform 0 1 1487 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_45
timestamp 1757161594
transform 0 1 2887 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_46
timestamp 1757161594
transform 0 1 3167 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_47
timestamp 1757161594
transform 0 1 2607 1 0 7838
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_0
timestamp 1757161594
transform 0 1 647 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_1
timestamp 1757161594
transform 0 1 927 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_2
timestamp 1757161594
transform 0 1 367 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_3
timestamp 1757161594
transform 0 1 87 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_4
timestamp 1757161594
transform 0 1 2047 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_5
timestamp 1757161594
transform 0 1 2327 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_6
timestamp 1757161594
transform 0 1 1767 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_7
timestamp 1757161594
transform 0 1 1207 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_8
timestamp 1757161594
transform 0 1 1487 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9
timestamp 1757161594
transform 0 1 367 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_10
timestamp 1757161594
transform 0 1 647 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_11
timestamp 1757161594
transform 0 1 927 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_12
timestamp 1757161594
transform 0 1 2887 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_13
timestamp 1757161594
transform 0 1 3167 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_14
timestamp 1757161594
transform 0 1 2607 1 0 9148
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_15
timestamp 1757161594
transform 0 1 87 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_16
timestamp 1757161594
transform 0 1 2047 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_17
timestamp 1757161594
transform 0 1 2327 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_18
timestamp 1757161594
transform 0 1 1767 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_19
timestamp 1757161594
transform 0 1 1207 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_20
timestamp 1757161594
transform 0 1 1487 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_21
timestamp 1757161594
transform 0 1 2607 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_22
timestamp 1757161594
transform 0 1 2887 1 0 -172
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGYFYD  sky130_fd_pr__nfet_01v8_lvt_QGYFYD_23
timestamp 1757161594
transform 0 1 3167 1 0 -172
box -134 -107 134 107
<< labels >>
flabel metal3 s 3690 2140 3790 2240 0 FreeSans 782 0 0 0 Vref
port 0 nsew
<< end >>
