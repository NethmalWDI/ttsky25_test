magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect 2020 730 13820 750
rect 2020 560 2120 730
rect 2160 560 13820 730
rect 2020 -720 13820 560
rect 2020 -920 7740 -720
rect 7860 -920 13820 -720
rect 2020 -1420 13820 -920
rect 2020 -1620 7720 -1420
rect 8200 -1620 13820 -1420
rect 2020 -2120 13820 -1620
rect 2020 -2320 7700 -2120
rect 8180 -2320 13820 -2120
rect 2020 -2740 13820 -2320
rect 2020 -2980 7740 -2740
rect 8060 -2980 13820 -2740
rect 2020 -3660 13820 -2980
rect 1870 -3840 13820 -3660
rect 1870 -4070 2130 -3840
rect 2150 -3850 2230 -3840
rect 6636 -3860 6724 -3840
rect 7820 -3850 7940 -3840
rect 13640 -3910 13820 -3840
<< pwell >>
rect 2014 -5146 2476 -5044
rect 2834 -8946 3056 -8264
<< psubdiff >>
rect 2040 -5120 2450 -5070
rect 2860 -8345 3030 -8290
rect 2860 -8379 2883 -8345
rect 2917 -8379 3030 -8345
rect 2860 -8413 3030 -8379
rect 2860 -8447 2883 -8413
rect 2917 -8447 3030 -8413
rect 2860 -8481 3030 -8447
rect 2860 -8515 2883 -8481
rect 2917 -8515 3030 -8481
rect 2860 -8549 3030 -8515
rect 2860 -8583 2883 -8549
rect 2917 -8583 3030 -8549
rect 2860 -8617 3030 -8583
rect 2860 -8651 2883 -8617
rect 2917 -8651 3030 -8617
rect 2860 -8685 3030 -8651
rect 2860 -8719 2883 -8685
rect 2917 -8719 3030 -8685
rect 2860 -8753 3030 -8719
rect 2860 -8787 2883 -8753
rect 2917 -8787 3030 -8753
rect 2860 -8821 3030 -8787
rect 2860 -8855 2883 -8821
rect 2917 -8855 3030 -8821
rect 2860 -8920 3030 -8855
<< nsubdiff >>
rect 10900 424 12000 480
rect 10900 322 10954 424
rect 11940 322 12000 424
rect 10900 300 12000 322
rect 7860 -3451 7910 -3390
rect 7860 -3485 7868 -3451
rect 7902 -3485 7910 -3451
rect 7860 -3519 7910 -3485
rect 7860 -3553 7868 -3519
rect 7902 -3553 7910 -3519
rect 7860 -3587 7910 -3553
rect 7860 -3621 7868 -3587
rect 7902 -3621 7910 -3587
rect 7860 -3655 7910 -3621
rect 7860 -3689 7868 -3655
rect 7902 -3689 7910 -3655
rect 7860 -3750 7910 -3689
<< psubdiffcont >>
rect 2883 -8379 2917 -8345
rect 2883 -8447 2917 -8413
rect 2883 -8515 2917 -8481
rect 2883 -8583 2917 -8549
rect 2883 -8651 2917 -8617
rect 2883 -8719 2917 -8685
rect 2883 -8787 2917 -8753
rect 2883 -8855 2917 -8821
<< nsubdiffcont >>
rect 10954 322 11940 424
rect 7868 -3485 7902 -3451
rect 7868 -3553 7902 -3519
rect 7868 -3621 7902 -3587
rect 7868 -3689 7902 -3655
<< locali >>
rect 7280 737 8980 750
rect 7280 710 7321 737
rect 6960 703 7321 710
rect 7355 703 7393 737
rect 7427 703 7465 737
rect 7499 703 7537 737
rect 7571 703 7609 737
rect 7643 703 7681 737
rect 7715 703 7753 737
rect 7787 703 7825 737
rect 7859 703 7897 737
rect 7931 703 7969 737
rect 8003 703 8041 737
rect 8075 703 8113 737
rect 8147 703 8185 737
rect 8219 703 8257 737
rect 8291 703 8329 737
rect 8363 703 8401 737
rect 8435 703 8473 737
rect 8507 703 8545 737
rect 8579 703 8617 737
rect 8651 703 8689 737
rect 8723 703 8761 737
rect 8795 703 8833 737
rect 8867 703 8905 737
rect 8939 710 8980 737
rect 8939 703 9620 710
rect 6960 680 9620 703
rect 10900 426 12000 480
rect 10900 424 10962 426
rect 11932 424 12000 426
rect 10900 322 10954 424
rect 11940 322 12000 424
rect 10900 320 10962 322
rect 11932 320 12000 322
rect 10900 300 12000 320
rect 13000 197 13540 200
rect 13000 163 13037 197
rect 13071 163 13109 197
rect 13143 163 13181 197
rect 13215 163 13253 197
rect 13287 163 13325 197
rect 13359 163 13397 197
rect 13431 163 13469 197
rect 13503 163 13540 197
rect 13000 150 13540 163
rect 7860 -3445 7910 -3390
rect 7860 -3485 7868 -3445
rect 7902 -3485 7910 -3445
rect 7860 -3517 7910 -3485
rect 7860 -3553 7868 -3517
rect 7902 -3553 7910 -3517
rect 7860 -3587 7910 -3553
rect 7860 -3623 7868 -3587
rect 7902 -3623 7910 -3587
rect 7860 -3655 7910 -3623
rect 7860 -3695 7868 -3655
rect 7902 -3695 7910 -3655
rect 7860 -3750 7910 -3695
rect 2020 -5076 2610 -5060
rect 2020 -5078 2497 -5076
rect 2020 -5112 2048 -5078
rect 2082 -5112 2120 -5078
rect 2154 -5112 2192 -5078
rect 2226 -5112 2264 -5078
rect 2298 -5112 2336 -5078
rect 2370 -5112 2408 -5078
rect 2442 -5110 2497 -5078
rect 2531 -5110 2610 -5076
rect 2442 -5112 2610 -5110
rect 2020 -5140 2610 -5112
rect 2860 -8296 3030 -8290
rect 2860 -8330 2993 -8296
rect 3027 -8330 3030 -8296
rect 2860 -8331 3030 -8330
rect 2860 -8379 2883 -8331
rect 2917 -8368 3030 -8331
rect 2917 -8379 2993 -8368
rect 2860 -8402 2993 -8379
rect 3027 -8402 3030 -8368
rect 2860 -8403 3030 -8402
rect 2860 -8447 2883 -8403
rect 2917 -8440 3030 -8403
rect 2917 -8447 2993 -8440
rect 2860 -8474 2993 -8447
rect 3027 -8474 3030 -8440
rect 2860 -8475 3030 -8474
rect 2860 -8515 2883 -8475
rect 2917 -8512 3030 -8475
rect 2917 -8515 2993 -8512
rect 2860 -8546 2993 -8515
rect 3027 -8546 3030 -8512
rect 2860 -8547 3030 -8546
rect 2860 -8583 2883 -8547
rect 2917 -8583 3030 -8547
rect 2860 -8584 3030 -8583
rect 2860 -8617 2993 -8584
rect 2860 -8653 2883 -8617
rect 2917 -8618 2993 -8617
rect 3027 -8618 3030 -8584
rect 2917 -8653 3030 -8618
rect 2860 -8656 3030 -8653
rect 2860 -8685 2993 -8656
rect 2860 -8725 2883 -8685
rect 2917 -8690 2993 -8685
rect 3027 -8690 3030 -8656
rect 2917 -8725 3030 -8690
rect 2860 -8728 3030 -8725
rect 2860 -8753 2993 -8728
rect 2860 -8797 2883 -8753
rect 2917 -8762 2993 -8753
rect 3027 -8762 3030 -8728
rect 2917 -8797 3030 -8762
rect 2860 -8800 3030 -8797
rect 2860 -8821 2993 -8800
rect 2860 -8869 2883 -8821
rect 2917 -8834 2993 -8821
rect 3027 -8834 3030 -8800
rect 2917 -8869 3030 -8834
rect 2860 -8920 3030 -8869
<< viali >>
rect 7321 703 7355 737
rect 7393 703 7427 737
rect 7465 703 7499 737
rect 7537 703 7571 737
rect 7609 703 7643 737
rect 7681 703 7715 737
rect 7753 703 7787 737
rect 7825 703 7859 737
rect 7897 703 7931 737
rect 7969 703 8003 737
rect 8041 703 8075 737
rect 8113 703 8147 737
rect 8185 703 8219 737
rect 8257 703 8291 737
rect 8329 703 8363 737
rect 8401 703 8435 737
rect 8473 703 8507 737
rect 8545 703 8579 737
rect 8617 703 8651 737
rect 8689 703 8723 737
rect 8761 703 8795 737
rect 8833 703 8867 737
rect 8905 703 8939 737
rect 10962 424 11932 426
rect 10962 322 11932 424
rect 10962 320 11932 322
rect 13037 163 13071 197
rect 13109 163 13143 197
rect 13181 163 13215 197
rect 13253 163 13287 197
rect 13325 163 13359 197
rect 13397 163 13431 197
rect 13469 163 13503 197
rect 7868 -3451 7902 -3445
rect 7868 -3479 7902 -3451
rect 7868 -3519 7902 -3517
rect 7868 -3551 7902 -3519
rect 7868 -3621 7902 -3589
rect 7868 -3623 7902 -3621
rect 7868 -3689 7902 -3661
rect 7868 -3695 7902 -3689
rect 2048 -5112 2082 -5078
rect 2120 -5112 2154 -5078
rect 2192 -5112 2226 -5078
rect 2264 -5112 2298 -5078
rect 2336 -5112 2370 -5078
rect 2408 -5112 2442 -5078
rect 2497 -5110 2531 -5076
rect 2993 -8330 3027 -8296
rect 2883 -8345 2917 -8331
rect 2883 -8365 2917 -8345
rect 2993 -8402 3027 -8368
rect 2883 -8413 2917 -8403
rect 2883 -8437 2917 -8413
rect 2993 -8474 3027 -8440
rect 2883 -8481 2917 -8475
rect 2883 -8509 2917 -8481
rect 2993 -8546 3027 -8512
rect 2883 -8549 2917 -8547
rect 2883 -8581 2917 -8549
rect 2993 -8618 3027 -8584
rect 2883 -8651 2917 -8619
rect 2883 -8653 2917 -8651
rect 2993 -8690 3027 -8656
rect 2883 -8719 2917 -8691
rect 2883 -8725 2917 -8719
rect 2993 -8762 3027 -8728
rect 2883 -8787 2917 -8763
rect 2883 -8797 2917 -8787
rect 2993 -8834 3027 -8800
rect 2883 -8855 2917 -8835
rect 2883 -8869 2917 -8855
<< metal1 >>
rect 7280 737 8980 750
rect 7280 710 7321 737
rect 2020 703 7321 710
rect 7355 703 7393 737
rect 7427 703 7465 737
rect 7499 703 7537 737
rect 7571 703 7609 737
rect 7643 703 7681 737
rect 7715 703 7753 737
rect 7787 703 7825 737
rect 7859 703 7897 737
rect 7931 703 7969 737
rect 8003 703 8041 737
rect 8075 703 8113 737
rect 8147 703 8185 737
rect 8219 703 8257 737
rect 8291 703 8329 737
rect 8363 703 8401 737
rect 8435 703 8473 737
rect 8507 703 8545 737
rect 8579 703 8617 737
rect 8651 703 8689 737
rect 8723 703 8761 737
rect 8795 703 8833 737
rect 8867 703 8905 737
rect 8939 710 8980 737
rect 8939 703 12000 710
rect 2020 630 12000 703
rect 2020 300 2100 630
rect 2140 400 2200 630
rect 6203 578 6299 581
rect 6203 410 6303 578
rect 1890 276 1990 300
rect 1890 224 1914 276
rect 1966 224 1990 276
rect 1780 -1727 1860 -1700
rect 1780 -1779 1793 -1727
rect 1845 -1779 1860 -1727
rect 1670 -2425 1750 -2400
rect 1670 -2477 1682 -2425
rect 1734 -2477 1750 -2425
rect 1670 -4433 1750 -2477
rect 1780 -4323 1860 -1779
rect 1780 -4375 1794 -4323
rect 1846 -4375 1860 -4323
rect 1780 -4390 1860 -4375
rect 1670 -4485 1681 -4433
rect 1733 -4485 1750 -4433
rect 1670 -4500 1750 -4485
rect 1890 -4740 1990 224
rect 2020 120 2120 300
rect 3493 281 3994 357
rect 6247 286 6303 410
rect 6399 411 6480 630
rect 10491 578 10587 585
rect 10491 414 10591 578
rect 6399 386 6456 411
rect 10528 381 10591 414
rect 3493 229 3628 281
rect 3680 229 3692 281
rect 3744 229 3756 281
rect 3808 229 3820 281
rect 3872 229 3994 281
rect 3493 200 3994 229
rect 6230 271 6303 286
rect 6230 219 6240 271
rect 6292 219 6303 271
rect 6230 204 6303 219
rect 6247 200 6303 204
rect 7703 281 8204 361
rect 7703 229 7824 281
rect 7876 229 7888 281
rect 7940 229 7952 281
rect 8004 229 8016 281
rect 8068 229 8204 281
rect 7703 200 8204 229
rect 10535 278 10591 381
rect 10900 480 12000 630
rect 10900 426 13540 480
rect 10900 320 10962 426
rect 11932 320 13540 426
rect 10900 300 13540 320
rect 10535 226 10539 278
rect 10535 200 10591 226
rect 13000 197 13540 300
rect 13000 163 13037 197
rect 13071 163 13109 197
rect 13143 163 13181 197
rect 13215 163 13253 197
rect 13287 163 13325 197
rect 13359 163 13397 197
rect 13431 163 13469 197
rect 13503 163 13540 197
rect 13000 150 13540 163
rect 2020 60 13520 120
rect 2020 -553 2120 60
rect 2660 -340 2780 60
rect 3920 -340 4020 60
rect 5180 -340 5280 60
rect 6460 -340 6540 60
rect 7700 -340 7800 60
rect 8980 -340 9080 60
rect 10220 -340 10320 60
rect 11480 -340 11600 60
rect 12760 -340 12860 60
rect 13420 -340 13520 60
rect 2260 -400 2780 -340
rect 2920 -400 4020 -340
rect 4200 -400 5280 -340
rect 5440 -400 6540 -340
rect 6700 -400 7800 -340
rect 7980 -400 9080 -340
rect 9220 -400 10320 -340
rect 10480 -400 11600 -340
rect 11760 -400 12860 -340
rect 13020 -400 13520 -340
rect 2020 -605 2043 -553
rect 2095 -605 2120 -553
rect 2720 -560 2780 -400
rect 2020 -1231 2120 -605
rect 2260 -620 2780 -560
rect 2920 -553 3940 -540
rect 2920 -605 2951 -553
rect 3003 -605 3015 -553
rect 3067 -605 3079 -553
rect 3131 -605 3143 -553
rect 3195 -605 3207 -553
rect 3259 -605 3271 -553
rect 3323 -605 3335 -553
rect 3387 -605 3399 -553
rect 3451 -605 3463 -553
rect 3515 -605 3527 -553
rect 3579 -605 3591 -553
rect 3643 -605 3655 -553
rect 3707 -605 3719 -553
rect 3771 -605 3783 -553
rect 3835 -605 3847 -553
rect 3899 -605 3940 -553
rect 2920 -620 3940 -605
rect 4181 -557 5188 -541
rect 4181 -609 4210 -557
rect 4262 -609 4274 -557
rect 4326 -609 4338 -557
rect 4390 -609 4402 -557
rect 4454 -609 4466 -557
rect 4518 -609 4530 -557
rect 4582 -609 4594 -557
rect 4646 -609 4658 -557
rect 4710 -609 4722 -557
rect 4774 -609 4786 -557
rect 4838 -609 4850 -557
rect 4902 -609 4914 -557
rect 4966 -609 4978 -557
rect 5030 -609 5042 -557
rect 5094 -609 5106 -557
rect 5158 -609 5188 -557
rect 4181 -619 5188 -609
rect 5439 -555 6444 -543
rect 5439 -607 5474 -555
rect 5526 -607 5538 -555
rect 5590 -607 5602 -555
rect 5654 -607 5666 -555
rect 5718 -607 5730 -555
rect 5782 -607 5794 -555
rect 5846 -607 5858 -555
rect 5910 -607 5922 -555
rect 5974 -607 5986 -555
rect 6038 -607 6050 -555
rect 6102 -607 6114 -555
rect 6166 -607 6178 -555
rect 6230 -607 6242 -555
rect 6294 -607 6306 -555
rect 6358 -607 6370 -555
rect 6422 -607 6444 -555
rect 2700 -1020 2780 -620
rect 3980 -740 4080 -620
rect 5240 -740 5340 -620
rect 5439 -622 6444 -607
rect 6703 -559 7719 -545
rect 6703 -611 6738 -559
rect 6790 -611 6802 -559
rect 6854 -611 6866 -559
rect 6918 -611 6930 -559
rect 6982 -611 6994 -559
rect 7046 -611 7058 -559
rect 7110 -611 7122 -559
rect 7174 -611 7186 -559
rect 7238 -611 7250 -559
rect 7302 -611 7314 -559
rect 7366 -611 7378 -559
rect 7430 -611 7442 -559
rect 7494 -611 7506 -559
rect 7558 -611 7570 -559
rect 7622 -611 7634 -559
rect 7686 -611 7719 -559
rect 6703 -620 7719 -611
rect 7976 -557 8959 -543
rect 7976 -609 7993 -557
rect 8045 -609 8057 -557
rect 8109 -609 8121 -557
rect 8173 -609 8185 -557
rect 8237 -609 8249 -557
rect 8301 -609 8313 -557
rect 8365 -609 8377 -557
rect 8429 -609 8441 -557
rect 8493 -609 8505 -557
rect 8557 -609 8569 -557
rect 8621 -609 8633 -557
rect 8685 -609 8697 -557
rect 8749 -609 8761 -557
rect 8813 -609 8825 -557
rect 8877 -609 8889 -557
rect 8941 -609 8959 -557
rect 3970 -762 4080 -740
rect 3970 -814 3994 -762
rect 4046 -814 4080 -762
rect 3970 -826 4080 -814
rect 3970 -878 3994 -826
rect 4046 -878 4080 -826
rect 3970 -900 4080 -878
rect 5230 -762 5340 -740
rect 5230 -814 5254 -762
rect 5306 -814 5340 -762
rect 5230 -826 5340 -814
rect 5230 -878 5254 -826
rect 5306 -878 5340 -826
rect 5230 -900 5340 -878
rect 3980 -1020 4080 -900
rect 5240 -1020 5340 -900
rect 6500 -708 6640 -620
rect 6500 -760 6564 -708
rect 6616 -760 6640 -708
rect 7760 -740 7860 -620
rect 7976 -623 8959 -609
rect 9235 -557 10239 -547
rect 9235 -609 9264 -557
rect 9316 -609 9328 -557
rect 9380 -609 9392 -557
rect 9444 -609 9456 -557
rect 9508 -609 9520 -557
rect 9572 -609 9584 -557
rect 9636 -609 9648 -557
rect 9700 -609 9712 -557
rect 9764 -609 9776 -557
rect 9828 -609 9840 -557
rect 9892 -609 9904 -557
rect 9956 -609 9968 -557
rect 10020 -609 10032 -557
rect 10084 -609 10096 -557
rect 10148 -609 10160 -557
rect 10212 -609 10239 -557
rect 9020 -740 9120 -620
rect 9235 -622 10239 -609
rect 10501 -560 11503 -540
rect 10501 -612 10527 -560
rect 10579 -612 10591 -560
rect 10643 -612 10655 -560
rect 10707 -612 10719 -560
rect 10771 -612 10783 -560
rect 10835 -612 10847 -560
rect 10899 -612 10911 -560
rect 10963 -612 10975 -560
rect 11027 -612 11039 -560
rect 11091 -612 11103 -560
rect 11155 -612 11167 -560
rect 11219 -612 11231 -560
rect 11283 -612 11295 -560
rect 11347 -612 11359 -560
rect 11411 -612 11423 -560
rect 11475 -612 11503 -560
rect 6500 -772 6640 -760
rect 6500 -824 6564 -772
rect 6616 -824 6640 -772
rect 6500 -836 6640 -824
rect 6500 -888 6564 -836
rect 6616 -888 6640 -836
rect 6500 -900 6640 -888
rect 7750 -762 7860 -740
rect 7750 -814 7774 -762
rect 7826 -814 7860 -762
rect 7750 -826 7860 -814
rect 7750 -878 7774 -826
rect 7826 -878 7860 -826
rect 7750 -900 7860 -878
rect 9010 -762 9120 -740
rect 9010 -814 9034 -762
rect 9086 -814 9120 -762
rect 9010 -826 9120 -814
rect 9010 -878 9034 -826
rect 9086 -878 9120 -826
rect 9010 -900 9120 -878
rect 6500 -952 6564 -900
rect 6616 -952 6640 -900
rect 6500 -1020 6640 -952
rect 7760 -1020 7860 -900
rect 9020 -1020 9120 -900
rect 10280 -724 10440 -620
rect 10501 -623 11503 -612
rect 11764 -560 12757 -538
rect 11764 -612 11790 -560
rect 11842 -612 11854 -560
rect 11906 -612 11918 -560
rect 11970 -612 11982 -560
rect 12034 -612 12046 -560
rect 12098 -612 12110 -560
rect 12162 -612 12174 -560
rect 12226 -612 12238 -560
rect 12290 -612 12302 -560
rect 12354 -612 12366 -560
rect 12418 -612 12430 -560
rect 12482 -612 12494 -560
rect 12546 -612 12558 -560
rect 12610 -612 12622 -560
rect 12674 -612 12686 -560
rect 12738 -612 12757 -560
rect 13460 -580 13520 -400
rect 10280 -776 10356 -724
rect 10408 -776 10440 -724
rect 10280 -788 10440 -776
rect 10280 -840 10356 -788
rect 10408 -840 10440 -788
rect 10280 -852 10440 -840
rect 10280 -904 10356 -852
rect 10408 -904 10440 -852
rect 10280 -916 10440 -904
rect 10280 -968 10356 -916
rect 10408 -968 10440 -916
rect 2150 -1048 2230 -1040
rect 2149 -1055 2230 -1048
rect 2149 -1107 2162 -1055
rect 2214 -1107 2230 -1055
rect 2280 -1080 2780 -1020
rect 2149 -1113 2230 -1107
rect 2020 -1283 2044 -1231
rect 2096 -1283 2120 -1231
rect 2020 -1915 2120 -1283
rect 2020 -1967 2044 -1915
rect 2096 -1967 2120 -1915
rect 2020 -2616 2120 -1967
rect 2020 -2668 2045 -2616
rect 2097 -2668 2120 -2616
rect 2020 -2680 2120 -2668
rect 2020 -3106 2100 -3080
rect 2020 -3158 2032 -3106
rect 2084 -3158 2100 -3106
rect 2020 -4546 2100 -3158
rect 2150 -4213 2230 -1113
rect 2720 -1240 2780 -1080
rect 2920 -1048 3920 -1040
rect 2920 -1100 2993 -1048
rect 3045 -1100 3057 -1048
rect 3109 -1100 3121 -1048
rect 3173 -1100 3185 -1048
rect 3237 -1100 3249 -1048
rect 3301 -1100 3313 -1048
rect 3365 -1100 3377 -1048
rect 3429 -1100 3441 -1048
rect 3493 -1100 3505 -1048
rect 3557 -1100 3569 -1048
rect 3621 -1100 3633 -1048
rect 3685 -1100 3697 -1048
rect 3749 -1100 3761 -1048
rect 3813 -1100 3825 -1048
rect 3877 -1100 3920 -1048
rect 2920 -1120 3920 -1100
rect 2280 -1320 2780 -1240
rect 2920 -1236 3940 -1220
rect 2920 -1288 2951 -1236
rect 3003 -1288 3015 -1236
rect 3067 -1288 3079 -1236
rect 3131 -1288 3143 -1236
rect 3195 -1288 3207 -1236
rect 3259 -1288 3271 -1236
rect 3323 -1288 3335 -1236
rect 3387 -1288 3399 -1236
rect 3451 -1288 3463 -1236
rect 3515 -1288 3527 -1236
rect 3579 -1288 3591 -1236
rect 3643 -1288 3655 -1236
rect 3707 -1288 3719 -1236
rect 3771 -1288 3783 -1236
rect 3835 -1288 3847 -1236
rect 3899 -1288 3940 -1236
rect 2920 -1300 3940 -1288
rect 4000 -1320 4080 -1020
rect 4180 -1050 5180 -1040
rect 4180 -1102 4239 -1050
rect 4291 -1102 4303 -1050
rect 4355 -1102 4367 -1050
rect 4419 -1102 4431 -1050
rect 4483 -1102 4495 -1050
rect 4547 -1102 4559 -1050
rect 4611 -1102 4623 -1050
rect 4675 -1102 4687 -1050
rect 4739 -1102 4751 -1050
rect 4803 -1102 4815 -1050
rect 4867 -1102 4879 -1050
rect 4931 -1102 4943 -1050
rect 4995 -1102 5007 -1050
rect 5059 -1102 5071 -1050
rect 5123 -1102 5180 -1050
rect 4180 -1120 5180 -1102
rect 5260 -1046 5340 -1020
rect 5460 -1037 6440 -1024
rect 5460 -1038 6448 -1037
rect 5260 -1054 5342 -1046
rect 5260 -1106 5275 -1054
rect 5327 -1106 5342 -1054
rect 5460 -1090 5481 -1038
rect 5533 -1090 5545 -1038
rect 5597 -1090 5609 -1038
rect 5661 -1090 5673 -1038
rect 5725 -1090 5737 -1038
rect 5789 -1090 5801 -1038
rect 5853 -1090 5865 -1038
rect 5917 -1090 5929 -1038
rect 5981 -1090 5993 -1038
rect 6045 -1090 6057 -1038
rect 6109 -1090 6121 -1038
rect 6173 -1090 6185 -1038
rect 6237 -1090 6249 -1038
rect 6301 -1090 6313 -1038
rect 6365 -1090 6377 -1038
rect 6429 -1090 6448 -1038
rect 5460 -1098 6440 -1090
rect 5260 -1114 5342 -1106
rect 4182 -1242 5183 -1218
rect 4182 -1294 4220 -1242
rect 4272 -1294 4284 -1242
rect 4336 -1294 4348 -1242
rect 4400 -1294 4412 -1242
rect 4464 -1294 4476 -1242
rect 4528 -1294 4540 -1242
rect 4592 -1294 4604 -1242
rect 4656 -1294 4668 -1242
rect 4720 -1294 4732 -1242
rect 4784 -1294 4796 -1242
rect 4848 -1294 4860 -1242
rect 4912 -1294 4924 -1242
rect 4976 -1294 4988 -1242
rect 5040 -1294 5052 -1242
rect 5104 -1294 5116 -1242
rect 5168 -1294 5183 -1242
rect 4182 -1311 5183 -1294
rect 5260 -1300 5340 -1114
rect 6520 -1140 6640 -1020
rect 6700 -1046 7680 -1040
rect 6700 -1098 6746 -1046
rect 6798 -1098 6810 -1046
rect 6862 -1098 6874 -1046
rect 6926 -1098 6938 -1046
rect 6990 -1098 7002 -1046
rect 7054 -1098 7066 -1046
rect 7118 -1098 7130 -1046
rect 7182 -1098 7194 -1046
rect 7246 -1098 7258 -1046
rect 7310 -1098 7322 -1046
rect 7374 -1098 7386 -1046
rect 7438 -1098 7450 -1046
rect 7502 -1098 7514 -1046
rect 7566 -1098 7578 -1046
rect 7630 -1098 7680 -1046
rect 6700 -1120 7680 -1098
rect 2700 -1700 2780 -1320
rect 3980 -1440 4080 -1320
rect 3970 -1462 4080 -1440
rect 3970 -1514 3994 -1462
rect 4046 -1514 4080 -1462
rect 3970 -1526 4080 -1514
rect 3970 -1578 3994 -1526
rect 4046 -1578 4080 -1526
rect 3970 -1600 4080 -1578
rect 2280 -1780 2780 -1700
rect 3980 -1720 4080 -1600
rect 5240 -1440 5340 -1300
rect 5460 -1237 6441 -1224
rect 5460 -1289 5498 -1237
rect 5550 -1289 5562 -1237
rect 5614 -1289 5626 -1237
rect 5678 -1289 5690 -1237
rect 5742 -1289 5754 -1237
rect 5806 -1289 5818 -1237
rect 5870 -1289 5882 -1237
rect 5934 -1289 5946 -1237
rect 5998 -1289 6010 -1237
rect 6062 -1289 6074 -1237
rect 6126 -1289 6138 -1237
rect 6190 -1289 6202 -1237
rect 6254 -1289 6266 -1237
rect 6318 -1289 6330 -1237
rect 6382 -1289 6441 -1237
rect 5460 -1309 6441 -1289
rect 6520 -1320 6600 -1140
rect 6700 -1237 7724 -1217
rect 6700 -1289 6737 -1237
rect 6789 -1289 6801 -1237
rect 6853 -1289 6865 -1237
rect 6917 -1289 6929 -1237
rect 6981 -1289 6993 -1237
rect 7045 -1289 7057 -1237
rect 7109 -1289 7121 -1237
rect 7173 -1289 7185 -1237
rect 7237 -1289 7249 -1237
rect 7301 -1289 7313 -1237
rect 7365 -1289 7377 -1237
rect 7429 -1289 7441 -1237
rect 7493 -1289 7505 -1237
rect 7557 -1289 7569 -1237
rect 7621 -1289 7633 -1237
rect 7685 -1289 7724 -1237
rect 6700 -1306 7724 -1289
rect 7780 -1300 7860 -1020
rect 7980 -1046 8960 -1040
rect 7980 -1098 8004 -1046
rect 8056 -1098 8068 -1046
rect 8120 -1098 8132 -1046
rect 8184 -1098 8196 -1046
rect 8248 -1098 8260 -1046
rect 8312 -1098 8324 -1046
rect 8376 -1098 8388 -1046
rect 8440 -1098 8452 -1046
rect 8504 -1098 8516 -1046
rect 8568 -1098 8580 -1046
rect 8632 -1098 8644 -1046
rect 8696 -1098 8708 -1046
rect 8760 -1098 8772 -1046
rect 8824 -1098 8836 -1046
rect 8888 -1098 8960 -1046
rect 7980 -1120 8960 -1098
rect 9040 -1054 9120 -1020
rect 9040 -1106 9053 -1054
rect 9105 -1106 9120 -1054
rect 9240 -1028 10240 -1020
rect 9240 -1034 10243 -1028
rect 9240 -1086 9267 -1034
rect 9319 -1086 9331 -1034
rect 9383 -1086 9395 -1034
rect 9447 -1086 9459 -1034
rect 9511 -1086 9523 -1034
rect 9575 -1086 9587 -1034
rect 9639 -1086 9651 -1034
rect 9703 -1086 9715 -1034
rect 9767 -1086 9779 -1034
rect 9831 -1086 9843 -1034
rect 9895 -1086 9907 -1034
rect 9959 -1086 9971 -1034
rect 10023 -1086 10035 -1034
rect 10087 -1086 10099 -1034
rect 10151 -1086 10163 -1034
rect 10215 -1086 10243 -1034
rect 10280 -1040 10440 -968
rect 11540 -740 11640 -620
rect 11764 -625 12757 -612
rect 12820 -740 12920 -620
rect 13040 -640 13520 -580
rect 11540 -762 11650 -740
rect 11540 -814 11574 -762
rect 11626 -814 11650 -762
rect 11540 -826 11650 -814
rect 11540 -878 11574 -826
rect 11626 -878 11650 -826
rect 11540 -900 11650 -878
rect 12810 -762 12920 -740
rect 12810 -814 12834 -762
rect 12886 -814 12920 -762
rect 12810 -826 12920 -814
rect 12810 -878 12834 -826
rect 12886 -878 12920 -826
rect 12810 -900 12920 -878
rect 11540 -1020 11640 -900
rect 12820 -1020 12920 -900
rect 9240 -1092 10243 -1086
rect 9240 -1100 10240 -1092
rect 6717 -1313 7723 -1306
rect 5240 -1462 5350 -1440
rect 5240 -1514 5274 -1462
rect 5326 -1514 5350 -1462
rect 5240 -1526 5350 -1514
rect 5240 -1578 5274 -1526
rect 5326 -1578 5350 -1526
rect 5240 -1600 5350 -1578
rect 5240 -1700 5340 -1600
rect 2720 -1940 2780 -1780
rect 2920 -1732 3920 -1720
rect 2920 -1784 2974 -1732
rect 3026 -1784 3038 -1732
rect 3090 -1784 3102 -1732
rect 3154 -1784 3166 -1732
rect 3218 -1784 3230 -1732
rect 3282 -1784 3294 -1732
rect 3346 -1784 3358 -1732
rect 3410 -1784 3422 -1732
rect 3474 -1784 3486 -1732
rect 3538 -1784 3550 -1732
rect 3602 -1784 3614 -1732
rect 3666 -1784 3678 -1732
rect 3730 -1784 3742 -1732
rect 3794 -1784 3806 -1732
rect 3858 -1784 3920 -1732
rect 2920 -1800 3920 -1784
rect 2280 -2000 2780 -1940
rect 2700 -2400 2780 -2000
rect 2920 -1911 3921 -1898
rect 2920 -1963 2950 -1911
rect 3002 -1963 3014 -1911
rect 3066 -1963 3078 -1911
rect 3130 -1963 3142 -1911
rect 3194 -1963 3206 -1911
rect 3258 -1963 3270 -1911
rect 3322 -1963 3334 -1911
rect 3386 -1963 3398 -1911
rect 3450 -1963 3462 -1911
rect 3514 -1963 3526 -1911
rect 3578 -1963 3590 -1911
rect 3642 -1963 3654 -1911
rect 3706 -1963 3718 -1911
rect 3770 -1963 3782 -1911
rect 3834 -1963 3846 -1911
rect 3898 -1963 3921 -1911
rect 2920 -2002 3921 -1963
rect 4000 -2000 4080 -1720
rect 4180 -1727 5180 -1720
rect 4180 -1779 4243 -1727
rect 4295 -1779 4307 -1727
rect 4359 -1779 4371 -1727
rect 4423 -1779 4435 -1727
rect 4487 -1779 4499 -1727
rect 4551 -1779 4563 -1727
rect 4615 -1779 4627 -1727
rect 4679 -1779 4691 -1727
rect 4743 -1779 4755 -1727
rect 4807 -1779 4819 -1727
rect 4871 -1779 4883 -1727
rect 4935 -1779 4947 -1727
rect 4999 -1779 5011 -1727
rect 5063 -1779 5075 -1727
rect 5127 -1779 5180 -1727
rect 4180 -1800 5180 -1779
rect 4180 -1921 5191 -1896
rect 4180 -1973 4216 -1921
rect 4268 -1973 4280 -1921
rect 4332 -1973 4344 -1921
rect 4396 -1973 4408 -1921
rect 4460 -1973 4472 -1921
rect 4524 -1973 4536 -1921
rect 4588 -1973 4600 -1921
rect 4652 -1973 4664 -1921
rect 4716 -1973 4728 -1921
rect 4780 -1973 4792 -1921
rect 4844 -1973 4856 -1921
rect 4908 -1973 4920 -1921
rect 4972 -1973 4984 -1921
rect 5036 -1973 5048 -1921
rect 5100 -1973 5112 -1921
rect 5164 -1973 5191 -1921
rect 4180 -1999 5191 -1973
rect 5260 -2000 5340 -1700
rect 5460 -1720 6436 -1718
rect 6500 -1720 6600 -1320
rect 7760 -1420 7860 -1300
rect 7985 -1231 8982 -1222
rect 7985 -1283 8020 -1231
rect 8072 -1283 8084 -1231
rect 8136 -1283 8148 -1231
rect 8200 -1283 8212 -1231
rect 8264 -1283 8276 -1231
rect 8328 -1283 8340 -1231
rect 8392 -1283 8404 -1231
rect 8456 -1283 8468 -1231
rect 8520 -1283 8532 -1231
rect 8584 -1283 8596 -1231
rect 8648 -1283 8660 -1231
rect 8712 -1283 8724 -1231
rect 8776 -1283 8788 -1231
rect 8840 -1283 8852 -1231
rect 8904 -1283 8982 -1231
rect 7985 -1311 8982 -1283
rect 9040 -1300 9120 -1106
rect 10300 -1140 10440 -1040
rect 10500 -1049 11500 -1020
rect 10500 -1101 10548 -1049
rect 10600 -1101 10612 -1049
rect 10664 -1101 10676 -1049
rect 10728 -1101 10740 -1049
rect 10792 -1101 10804 -1049
rect 10856 -1101 10868 -1049
rect 10920 -1101 10932 -1049
rect 10984 -1101 10996 -1049
rect 11048 -1101 11060 -1049
rect 11112 -1101 11124 -1049
rect 11176 -1101 11188 -1049
rect 11240 -1101 11252 -1049
rect 11304 -1101 11316 -1049
rect 11368 -1101 11380 -1049
rect 11432 -1101 11500 -1049
rect 10500 -1120 11500 -1101
rect 9020 -1440 9120 -1300
rect 9242 -1243 10232 -1222
rect 9242 -1295 9283 -1243
rect 9335 -1295 9347 -1243
rect 9399 -1295 9411 -1243
rect 9463 -1295 9475 -1243
rect 9527 -1295 9539 -1243
rect 9591 -1295 9603 -1243
rect 9655 -1295 9667 -1243
rect 9719 -1295 9731 -1243
rect 9783 -1295 9795 -1243
rect 9847 -1295 9859 -1243
rect 9911 -1295 9923 -1243
rect 9975 -1295 9987 -1243
rect 10039 -1295 10051 -1243
rect 10103 -1295 10115 -1243
rect 10167 -1295 10232 -1243
rect 9242 -1304 10232 -1295
rect 10300 -1300 10380 -1140
rect 9020 -1462 9130 -1440
rect 9020 -1514 9054 -1462
rect 9106 -1514 9130 -1462
rect 9020 -1526 9130 -1514
rect 9020 -1578 9054 -1526
rect 9106 -1578 9130 -1526
rect 9020 -1600 9130 -1578
rect 7760 -1700 7860 -1620
rect 9020 -1700 9120 -1600
rect 10280 -1700 10380 -1300
rect 10503 -1243 11494 -1219
rect 10503 -1295 10525 -1243
rect 10577 -1295 10589 -1243
rect 10641 -1295 10653 -1243
rect 10705 -1295 10717 -1243
rect 10769 -1295 10781 -1243
rect 10833 -1295 10845 -1243
rect 10897 -1295 10909 -1243
rect 10961 -1295 10973 -1243
rect 11025 -1295 11037 -1243
rect 11089 -1295 11101 -1243
rect 11153 -1295 11165 -1243
rect 11217 -1295 11229 -1243
rect 11281 -1295 11293 -1243
rect 11345 -1295 11357 -1243
rect 11409 -1295 11421 -1243
rect 11473 -1295 11494 -1243
rect 10503 -1316 11494 -1295
rect 11560 -1300 11640 -1020
rect 11760 -1056 12760 -1020
rect 11760 -1108 11814 -1056
rect 11866 -1108 11878 -1056
rect 11930 -1108 11942 -1056
rect 11994 -1108 12006 -1056
rect 12058 -1108 12070 -1056
rect 12122 -1108 12134 -1056
rect 12186 -1108 12198 -1056
rect 12250 -1108 12262 -1056
rect 12314 -1108 12326 -1056
rect 12378 -1108 12390 -1056
rect 12442 -1108 12454 -1056
rect 12506 -1108 12518 -1056
rect 12570 -1108 12582 -1056
rect 12634 -1108 12646 -1056
rect 12698 -1108 12760 -1056
rect 11760 -1120 12760 -1108
rect 11540 -1440 11640 -1300
rect 11757 -1237 12760 -1221
rect 11757 -1289 11783 -1237
rect 11835 -1289 11847 -1237
rect 11899 -1289 11911 -1237
rect 11963 -1289 11975 -1237
rect 12027 -1289 12039 -1237
rect 12091 -1289 12103 -1237
rect 12155 -1289 12167 -1237
rect 12219 -1289 12231 -1237
rect 12283 -1289 12295 -1237
rect 12347 -1289 12359 -1237
rect 12411 -1289 12423 -1237
rect 12475 -1289 12487 -1237
rect 12539 -1289 12551 -1237
rect 12603 -1289 12615 -1237
rect 12667 -1289 12679 -1237
rect 12731 -1289 12760 -1237
rect 11757 -1313 12760 -1289
rect 12840 -1300 12920 -1020
rect 13420 -1040 13520 -640
rect 13040 -1120 13520 -1040
rect 13460 -1260 13520 -1120
rect 12820 -1440 12920 -1300
rect 13040 -1320 13520 -1260
rect 11540 -1462 11650 -1440
rect 11540 -1514 11574 -1462
rect 11626 -1514 11650 -1462
rect 11540 -1526 11650 -1514
rect 11540 -1578 11574 -1526
rect 11626 -1578 11650 -1526
rect 11540 -1600 11650 -1578
rect 12810 -1462 12920 -1440
rect 12810 -1514 12834 -1462
rect 12886 -1514 12920 -1462
rect 12810 -1526 12920 -1514
rect 12810 -1578 12834 -1526
rect 12886 -1578 12920 -1526
rect 12810 -1600 12920 -1578
rect 11540 -1700 11640 -1600
rect 12820 -1700 12920 -1600
rect 5460 -1760 6460 -1720
rect 6520 -1760 6600 -1720
rect 5460 -1800 6600 -1760
rect 6720 -1737 7700 -1720
rect 6720 -1789 6762 -1737
rect 6814 -1789 6826 -1737
rect 6878 -1789 6890 -1737
rect 6942 -1789 6954 -1737
rect 7006 -1789 7018 -1737
rect 7070 -1789 7082 -1737
rect 7134 -1789 7146 -1737
rect 7198 -1789 7210 -1737
rect 7262 -1789 7274 -1737
rect 7326 -1789 7338 -1737
rect 7390 -1789 7402 -1737
rect 7454 -1789 7466 -1737
rect 7518 -1789 7530 -1737
rect 7582 -1789 7594 -1737
rect 7646 -1789 7700 -1737
rect 6720 -1800 7700 -1789
rect 5440 -1913 6460 -1901
rect 5440 -1965 5480 -1913
rect 5532 -1965 5544 -1913
rect 5596 -1965 5608 -1913
rect 5660 -1965 5672 -1913
rect 5724 -1965 5736 -1913
rect 5788 -1965 5800 -1913
rect 5852 -1965 5864 -1913
rect 5916 -1965 5928 -1913
rect 5980 -1965 5992 -1913
rect 6044 -1965 6056 -1913
rect 6108 -1965 6120 -1913
rect 6172 -1965 6184 -1913
rect 6236 -1965 6248 -1913
rect 6300 -1965 6312 -1913
rect 6364 -1965 6376 -1913
rect 6428 -1965 6460 -1913
rect 5440 -1999 6460 -1965
rect 6520 -2000 6600 -1800
rect 6711 -1922 7722 -1899
rect 6711 -1974 6739 -1922
rect 6791 -1974 6803 -1922
rect 6855 -1974 6867 -1922
rect 6919 -1974 6931 -1922
rect 6983 -1974 6995 -1922
rect 7047 -1974 7059 -1922
rect 7111 -1974 7123 -1922
rect 7175 -1974 7187 -1922
rect 7239 -1974 7251 -1922
rect 7303 -1974 7315 -1922
rect 7367 -1974 7379 -1922
rect 7431 -1974 7443 -1922
rect 7495 -1974 7507 -1922
rect 7559 -1974 7571 -1922
rect 7623 -1974 7635 -1922
rect 7687 -1974 7722 -1922
rect 6711 -1998 7722 -1974
rect 7780 -2000 7860 -1700
rect 7980 -1734 8960 -1720
rect 7980 -1786 8021 -1734
rect 8073 -1786 8085 -1734
rect 8137 -1786 8149 -1734
rect 8201 -1786 8213 -1734
rect 8265 -1786 8277 -1734
rect 8329 -1786 8341 -1734
rect 8393 -1786 8405 -1734
rect 8457 -1786 8469 -1734
rect 8521 -1786 8533 -1734
rect 8585 -1786 8597 -1734
rect 8649 -1786 8661 -1734
rect 8713 -1786 8725 -1734
rect 8777 -1786 8789 -1734
rect 8841 -1786 8853 -1734
rect 8905 -1786 8960 -1734
rect 7980 -1800 8960 -1786
rect 7970 -1923 8981 -1903
rect 7970 -1975 8000 -1923
rect 8052 -1975 8064 -1923
rect 8116 -1975 8128 -1923
rect 8180 -1975 8192 -1923
rect 8244 -1975 8256 -1923
rect 8308 -1975 8320 -1923
rect 8372 -1975 8384 -1923
rect 8436 -1975 8448 -1923
rect 8500 -1975 8512 -1923
rect 8564 -1975 8576 -1923
rect 8628 -1975 8640 -1923
rect 8692 -1975 8704 -1923
rect 8756 -1975 8768 -1923
rect 8820 -1975 8832 -1923
rect 8884 -1975 8896 -1923
rect 8948 -1975 8981 -1923
rect 7970 -1990 8981 -1975
rect 9040 -2000 9120 -1700
rect 9240 -1760 10240 -1720
rect 10300 -1760 10380 -1700
rect 9240 -1800 10380 -1760
rect 10500 -1727 11500 -1700
rect 10500 -1779 10566 -1727
rect 10618 -1779 10630 -1727
rect 10682 -1779 10694 -1727
rect 10746 -1779 10758 -1727
rect 10810 -1779 10822 -1727
rect 10874 -1779 10886 -1727
rect 10938 -1779 10950 -1727
rect 11002 -1779 11014 -1727
rect 11066 -1779 11078 -1727
rect 11130 -1779 11142 -1727
rect 11194 -1779 11206 -1727
rect 11258 -1779 11270 -1727
rect 11322 -1779 11334 -1727
rect 11386 -1779 11398 -1727
rect 11450 -1779 11500 -1727
rect 10500 -1800 11500 -1779
rect 9238 -1920 10240 -1905
rect 9238 -1972 9259 -1920
rect 9311 -1972 9323 -1920
rect 9375 -1972 9387 -1920
rect 9439 -1972 9451 -1920
rect 9503 -1972 9515 -1920
rect 9567 -1972 9579 -1920
rect 9631 -1972 9643 -1920
rect 9695 -1972 9707 -1920
rect 9759 -1972 9771 -1920
rect 9823 -1972 9835 -1920
rect 9887 -1972 9899 -1920
rect 9951 -1972 9963 -1920
rect 10015 -1972 10027 -1920
rect 10079 -1972 10091 -1920
rect 10143 -1972 10155 -1920
rect 10207 -1972 10240 -1920
rect 9238 -1989 10240 -1972
rect 10300 -2000 10380 -1800
rect 10497 -1924 11496 -1902
rect 10497 -1976 10521 -1924
rect 10573 -1976 10585 -1924
rect 10637 -1976 10649 -1924
rect 10701 -1976 10713 -1924
rect 10765 -1976 10777 -1924
rect 10829 -1976 10841 -1924
rect 10893 -1976 10905 -1924
rect 10957 -1976 10969 -1924
rect 11021 -1976 11033 -1924
rect 11085 -1976 11097 -1924
rect 11149 -1976 11161 -1924
rect 11213 -1976 11225 -1924
rect 11277 -1976 11289 -1924
rect 11341 -1976 11353 -1924
rect 11405 -1976 11417 -1924
rect 11469 -1976 11496 -1924
rect 10497 -1999 11496 -1976
rect 11560 -2000 11640 -1700
rect 11760 -1732 12760 -1700
rect 11760 -1784 11812 -1732
rect 11864 -1784 11876 -1732
rect 11928 -1784 11940 -1732
rect 11992 -1784 12004 -1732
rect 12056 -1784 12068 -1732
rect 12120 -1784 12132 -1732
rect 12184 -1784 12196 -1732
rect 12248 -1784 12260 -1732
rect 12312 -1784 12324 -1732
rect 12376 -1784 12388 -1732
rect 12440 -1784 12452 -1732
rect 12504 -1784 12516 -1732
rect 12568 -1784 12580 -1732
rect 12632 -1784 12644 -1732
rect 12696 -1784 12760 -1732
rect 11760 -1800 12760 -1784
rect 11762 -1921 12758 -1902
rect 11762 -1973 11780 -1921
rect 11832 -1973 11844 -1921
rect 11896 -1973 11908 -1921
rect 11960 -1973 11972 -1921
rect 12024 -1973 12036 -1921
rect 12088 -1973 12100 -1921
rect 12152 -1973 12164 -1921
rect 12216 -1973 12228 -1921
rect 12280 -1973 12292 -1921
rect 12344 -1973 12356 -1921
rect 12408 -1973 12420 -1921
rect 12472 -1973 12484 -1921
rect 12536 -1973 12548 -1921
rect 12600 -1973 12612 -1921
rect 12664 -1973 12676 -1921
rect 12728 -1973 12758 -1921
rect 11762 -1996 12758 -1973
rect 12840 -2000 12920 -1700
rect 13420 -1720 13520 -1320
rect 13880 -1052 13960 -1020
rect 13880 -1104 13892 -1052
rect 13944 -1104 13960 -1052
rect 13040 -1780 13520 -1720
rect 13460 -1940 13520 -1780
rect 13770 -1726 13850 -1700
rect 13770 -1778 13782 -1726
rect 13834 -1778 13850 -1726
rect 13040 -2000 13540 -1940
rect 3980 -2140 4080 -2000
rect 5240 -2140 5340 -2000
rect 3970 -2162 4080 -2140
rect 3970 -2214 3994 -2162
rect 4046 -2214 4080 -2162
rect 3970 -2226 4080 -2214
rect 3970 -2278 3994 -2226
rect 4046 -2278 4080 -2226
rect 3970 -2300 4080 -2278
rect 5230 -2162 5340 -2140
rect 5230 -2214 5254 -2162
rect 5306 -2214 5340 -2162
rect 5230 -2226 5340 -2214
rect 5230 -2278 5254 -2226
rect 5306 -2278 5340 -2226
rect 5230 -2300 5340 -2278
rect 3980 -2400 4080 -2300
rect 5240 -2400 5340 -2300
rect 6500 -2400 6600 -2000
rect 7760 -2120 7860 -2000
rect 9020 -2140 9120 -2000
rect 9020 -2162 9130 -2140
rect 9020 -2214 9054 -2162
rect 9106 -2214 9130 -2162
rect 9020 -2226 9130 -2214
rect 9020 -2278 9054 -2226
rect 9106 -2278 9130 -2226
rect 9020 -2300 9130 -2278
rect 7760 -2400 7860 -2320
rect 9020 -2400 9120 -2300
rect 10280 -2400 10380 -2000
rect 11540 -2140 11640 -2000
rect 12820 -2140 12920 -2000
rect 11540 -2162 11650 -2140
rect 11540 -2214 11574 -2162
rect 11626 -2214 11650 -2162
rect 11540 -2226 11650 -2214
rect 11540 -2278 11574 -2226
rect 11626 -2278 11650 -2226
rect 11540 -2300 11650 -2278
rect 12810 -2162 12920 -2140
rect 12810 -2214 12834 -2162
rect 12886 -2214 12920 -2162
rect 12810 -2226 12920 -2214
rect 12810 -2278 12834 -2226
rect 12886 -2278 12920 -2226
rect 12810 -2300 12920 -2278
rect 11540 -2400 11640 -2300
rect 12820 -2400 12920 -2300
rect 13460 -2400 13540 -2000
rect 2280 -2460 2780 -2400
rect 2720 -2620 2780 -2460
rect 2920 -2425 3920 -2400
rect 2920 -2477 2974 -2425
rect 3026 -2477 3038 -2425
rect 3090 -2477 3102 -2425
rect 3154 -2477 3166 -2425
rect 3218 -2477 3230 -2425
rect 3282 -2477 3294 -2425
rect 3346 -2477 3358 -2425
rect 3410 -2477 3422 -2425
rect 3474 -2477 3486 -2425
rect 3538 -2477 3550 -2425
rect 3602 -2477 3614 -2425
rect 3666 -2477 3678 -2425
rect 3730 -2477 3742 -2425
rect 3794 -2477 3806 -2425
rect 3858 -2477 3920 -2425
rect 2920 -2500 3920 -2477
rect 2280 -2680 2780 -2620
rect 2914 -2612 3925 -2603
rect 2914 -2664 2947 -2612
rect 2999 -2664 3011 -2612
rect 3063 -2664 3075 -2612
rect 3127 -2664 3139 -2612
rect 3191 -2664 3203 -2612
rect 3255 -2664 3267 -2612
rect 3319 -2664 3331 -2612
rect 3383 -2664 3395 -2612
rect 3447 -2664 3459 -2612
rect 3511 -2664 3523 -2612
rect 3575 -2664 3587 -2612
rect 3639 -2664 3651 -2612
rect 3703 -2664 3715 -2612
rect 3767 -2664 3779 -2612
rect 3831 -2664 3843 -2612
rect 3895 -2664 3925 -2612
rect 2914 -2679 3925 -2664
rect 4000 -2680 4080 -2400
rect 4179 -2420 5178 -2410
rect 4179 -2472 4250 -2420
rect 4302 -2472 4314 -2420
rect 4366 -2472 4378 -2420
rect 4430 -2472 4442 -2420
rect 4494 -2472 4506 -2420
rect 4558 -2472 4570 -2420
rect 4622 -2472 4634 -2420
rect 4686 -2472 4698 -2420
rect 4750 -2472 4762 -2420
rect 4814 -2472 4826 -2420
rect 4878 -2472 4890 -2420
rect 4942 -2472 4954 -2420
rect 5006 -2472 5018 -2420
rect 5070 -2472 5082 -2420
rect 5134 -2472 5178 -2420
rect 4179 -2509 5178 -2472
rect 2700 -3080 2780 -2680
rect 3980 -2800 4080 -2680
rect 4183 -2620 5199 -2603
rect 4183 -2672 4213 -2620
rect 4265 -2672 4277 -2620
rect 4329 -2672 4341 -2620
rect 4393 -2672 4405 -2620
rect 4457 -2672 4469 -2620
rect 4521 -2672 4533 -2620
rect 4585 -2672 4597 -2620
rect 4649 -2672 4661 -2620
rect 4713 -2672 4725 -2620
rect 4777 -2672 4789 -2620
rect 4841 -2672 4853 -2620
rect 4905 -2672 4917 -2620
rect 4969 -2672 4981 -2620
rect 5033 -2672 5045 -2620
rect 5097 -2672 5109 -2620
rect 5161 -2672 5199 -2620
rect 4183 -2683 5199 -2672
rect 5260 -2680 5340 -2400
rect 5460 -2440 6440 -2400
rect 6520 -2440 6600 -2400
rect 5460 -2480 6600 -2440
rect 6720 -2415 7700 -2400
rect 6720 -2467 6759 -2415
rect 6811 -2467 6823 -2415
rect 6875 -2467 6887 -2415
rect 6939 -2467 6951 -2415
rect 7003 -2467 7015 -2415
rect 7067 -2467 7079 -2415
rect 7131 -2467 7143 -2415
rect 7195 -2467 7207 -2415
rect 7259 -2467 7271 -2415
rect 7323 -2467 7335 -2415
rect 7387 -2467 7399 -2415
rect 7451 -2467 7463 -2415
rect 7515 -2467 7527 -2415
rect 7579 -2467 7591 -2415
rect 7643 -2467 7700 -2415
rect 6720 -2480 7700 -2467
rect 5437 -2620 6460 -2601
rect 5437 -2672 5479 -2620
rect 5531 -2672 5543 -2620
rect 5595 -2672 5607 -2620
rect 5659 -2672 5671 -2620
rect 5723 -2672 5735 -2620
rect 5787 -2672 5799 -2620
rect 5851 -2672 5863 -2620
rect 5915 -2672 5927 -2620
rect 5979 -2672 5991 -2620
rect 6043 -2672 6055 -2620
rect 6107 -2672 6119 -2620
rect 6171 -2672 6183 -2620
rect 6235 -2672 6247 -2620
rect 6299 -2672 6311 -2620
rect 6363 -2672 6375 -2620
rect 6427 -2672 6460 -2620
rect 5437 -2680 6460 -2672
rect 6520 -2680 6600 -2480
rect 6700 -2620 7719 -2603
rect 6700 -2672 6736 -2620
rect 6788 -2672 6800 -2620
rect 6852 -2672 6864 -2620
rect 6916 -2672 6928 -2620
rect 6980 -2672 6992 -2620
rect 7044 -2672 7056 -2620
rect 7108 -2672 7120 -2620
rect 7172 -2672 7184 -2620
rect 7236 -2672 7248 -2620
rect 7300 -2672 7312 -2620
rect 7364 -2672 7376 -2620
rect 7428 -2672 7440 -2620
rect 7492 -2672 7504 -2620
rect 7556 -2672 7568 -2620
rect 7620 -2672 7632 -2620
rect 7684 -2672 7719 -2620
rect 6700 -2680 7719 -2672
rect 7780 -2680 7860 -2400
rect 7980 -2406 8960 -2400
rect 7980 -2458 8009 -2406
rect 8061 -2458 8073 -2406
rect 8125 -2458 8137 -2406
rect 8189 -2458 8201 -2406
rect 8253 -2458 8265 -2406
rect 8317 -2458 8329 -2406
rect 8381 -2458 8393 -2406
rect 8445 -2458 8457 -2406
rect 8509 -2458 8521 -2406
rect 8573 -2458 8585 -2406
rect 8637 -2458 8649 -2406
rect 8701 -2458 8713 -2406
rect 8765 -2458 8777 -2406
rect 8829 -2458 8841 -2406
rect 8893 -2458 8960 -2406
rect 7980 -2480 8960 -2458
rect 5240 -2800 5340 -2680
rect 3970 -2822 4080 -2800
rect 3970 -2874 3994 -2822
rect 4046 -2874 4080 -2822
rect 3970 -2886 4080 -2874
rect 3970 -2938 3994 -2886
rect 4046 -2938 4080 -2886
rect 3970 -2960 4080 -2938
rect 5230 -2822 5340 -2800
rect 5230 -2874 5254 -2822
rect 5306 -2874 5340 -2822
rect 5230 -2886 5340 -2874
rect 5230 -2938 5254 -2886
rect 5306 -2938 5340 -2886
rect 5230 -2960 5340 -2938
rect 3980 -3080 4080 -2960
rect 5240 -3080 5340 -2960
rect 6500 -3080 6600 -2680
rect 7760 -2740 7860 -2680
rect 7977 -2620 8984 -2602
rect 7977 -2672 8004 -2620
rect 8056 -2672 8068 -2620
rect 8120 -2672 8132 -2620
rect 8184 -2672 8196 -2620
rect 8248 -2672 8260 -2620
rect 8312 -2672 8324 -2620
rect 8376 -2672 8388 -2620
rect 8440 -2672 8452 -2620
rect 8504 -2672 8516 -2620
rect 8568 -2672 8580 -2620
rect 8632 -2672 8644 -2620
rect 8696 -2672 8708 -2620
rect 8760 -2672 8772 -2620
rect 8824 -2672 8836 -2620
rect 8888 -2672 8900 -2620
rect 8952 -2672 8984 -2620
rect 7977 -2682 8984 -2672
rect 9040 -2680 9120 -2400
rect 9240 -2440 10240 -2400
rect 10300 -2440 10380 -2400
rect 9240 -2480 10380 -2440
rect 9020 -2800 9120 -2680
rect 9240 -2617 10240 -2604
rect 9240 -2669 9264 -2617
rect 9316 -2669 9328 -2617
rect 9380 -2669 9392 -2617
rect 9444 -2669 9456 -2617
rect 9508 -2669 9520 -2617
rect 9572 -2669 9584 -2617
rect 9636 -2669 9648 -2617
rect 9700 -2669 9712 -2617
rect 9764 -2669 9776 -2617
rect 9828 -2669 9840 -2617
rect 9892 -2669 9904 -2617
rect 9956 -2669 9968 -2617
rect 10020 -2669 10032 -2617
rect 10084 -2669 10096 -2617
rect 10148 -2669 10160 -2617
rect 10212 -2669 10240 -2617
rect 9240 -2681 10240 -2669
rect 10300 -2680 10380 -2480
rect 10500 -2424 11500 -2400
rect 10500 -2476 10564 -2424
rect 10616 -2476 10628 -2424
rect 10680 -2476 10692 -2424
rect 10744 -2476 10756 -2424
rect 10808 -2476 10820 -2424
rect 10872 -2476 10884 -2424
rect 10936 -2476 10948 -2424
rect 11000 -2476 11012 -2424
rect 11064 -2476 11076 -2424
rect 11128 -2476 11140 -2424
rect 11192 -2476 11204 -2424
rect 11256 -2476 11268 -2424
rect 11320 -2476 11332 -2424
rect 11384 -2476 11396 -2424
rect 11448 -2476 11500 -2424
rect 10500 -2500 11500 -2476
rect 9020 -2822 9130 -2800
rect 9020 -2874 9054 -2822
rect 9106 -2874 9130 -2822
rect 9020 -2886 9130 -2874
rect 9020 -2938 9054 -2886
rect 9106 -2938 9130 -2886
rect 9020 -2960 9130 -2938
rect 7760 -3080 7860 -2980
rect 9020 -3080 9120 -2960
rect 10280 -3060 10380 -2680
rect 10498 -2616 11499 -2598
rect 10498 -2668 10525 -2616
rect 10577 -2668 10589 -2616
rect 10641 -2668 10653 -2616
rect 10705 -2668 10717 -2616
rect 10769 -2668 10781 -2616
rect 10833 -2668 10845 -2616
rect 10897 -2668 10909 -2616
rect 10961 -2668 10973 -2616
rect 11025 -2668 11037 -2616
rect 11089 -2668 11101 -2616
rect 11153 -2668 11165 -2616
rect 11217 -2668 11229 -2616
rect 11281 -2668 11293 -2616
rect 11345 -2668 11357 -2616
rect 11409 -2668 11421 -2616
rect 11473 -2668 11499 -2616
rect 10498 -2682 11499 -2668
rect 11560 -2680 11640 -2400
rect 11760 -2429 12760 -2400
rect 11760 -2481 11812 -2429
rect 11864 -2481 11876 -2429
rect 11928 -2481 11940 -2429
rect 11992 -2481 12004 -2429
rect 12056 -2481 12068 -2429
rect 12120 -2481 12132 -2429
rect 12184 -2481 12196 -2429
rect 12248 -2481 12260 -2429
rect 12312 -2481 12324 -2429
rect 12376 -2481 12388 -2429
rect 12440 -2481 12452 -2429
rect 12504 -2481 12516 -2429
rect 12568 -2481 12580 -2429
rect 12632 -2481 12644 -2429
rect 12696 -2481 12760 -2429
rect 11760 -2500 12760 -2481
rect 2280 -3140 2780 -3080
rect 2720 -3300 2780 -3140
rect 2920 -3108 3920 -3080
rect 2920 -3160 2969 -3108
rect 3021 -3160 3033 -3108
rect 3085 -3160 3097 -3108
rect 3149 -3160 3161 -3108
rect 3213 -3160 3225 -3108
rect 3277 -3160 3289 -3108
rect 3341 -3160 3353 -3108
rect 3405 -3160 3417 -3108
rect 3469 -3160 3481 -3108
rect 3533 -3160 3545 -3108
rect 3597 -3160 3609 -3108
rect 3661 -3160 3673 -3108
rect 3725 -3160 3737 -3108
rect 3789 -3160 3801 -3108
rect 3853 -3160 3920 -3108
rect 2920 -3180 3920 -3160
rect 4000 -3227 4080 -3080
rect 4179 -3115 5182 -3091
rect 5260 -3112 5340 -3080
rect 4179 -3167 4248 -3115
rect 4300 -3167 4312 -3115
rect 4364 -3167 4376 -3115
rect 4428 -3167 4440 -3115
rect 4492 -3167 4504 -3115
rect 4556 -3167 4568 -3115
rect 4620 -3167 4632 -3115
rect 4684 -3167 4696 -3115
rect 4748 -3167 4760 -3115
rect 4812 -3167 4824 -3115
rect 4876 -3167 4888 -3115
rect 4940 -3167 4952 -3115
rect 5004 -3167 5016 -3115
rect 5068 -3167 5080 -3115
rect 5132 -3167 5182 -3115
rect 4179 -3180 5182 -3167
rect 5259 -3117 5340 -3112
rect 5259 -3169 5273 -3117
rect 5325 -3169 5340 -3117
rect 5444 -3096 6459 -3080
rect 5444 -3148 5474 -3096
rect 5526 -3148 5538 -3096
rect 5590 -3148 5602 -3096
rect 5654 -3148 5666 -3096
rect 5718 -3148 5730 -3096
rect 5782 -3148 5794 -3096
rect 5846 -3148 5858 -3096
rect 5910 -3148 5922 -3096
rect 5974 -3148 5986 -3096
rect 6038 -3148 6050 -3096
rect 6102 -3148 6114 -3096
rect 6166 -3148 6178 -3096
rect 6230 -3148 6242 -3096
rect 6294 -3148 6306 -3096
rect 6358 -3148 6370 -3096
rect 6422 -3148 6459 -3096
rect 5444 -3164 6459 -3148
rect 6720 -3104 7700 -3080
rect 6720 -3156 6726 -3104
rect 6778 -3156 6790 -3104
rect 6842 -3156 6854 -3104
rect 6906 -3156 6918 -3104
rect 6970 -3156 6982 -3104
rect 7034 -3156 7046 -3104
rect 7098 -3156 7110 -3104
rect 7162 -3156 7174 -3104
rect 7226 -3156 7238 -3104
rect 7290 -3156 7302 -3104
rect 7354 -3156 7366 -3104
rect 7418 -3156 7430 -3104
rect 7482 -3156 7494 -3104
rect 7546 -3156 7558 -3104
rect 7610 -3156 7622 -3104
rect 7674 -3156 7700 -3104
rect 5259 -3173 5340 -3169
rect 5260 -3224 5340 -3173
rect 6720 -3180 7700 -3156
rect 7780 -3246 7860 -3080
rect 7980 -3104 8960 -3080
rect 7980 -3156 7986 -3104
rect 8038 -3156 8050 -3104
rect 8102 -3156 8114 -3104
rect 8166 -3156 8178 -3104
rect 8230 -3156 8242 -3104
rect 8294 -3156 8306 -3104
rect 8358 -3156 8370 -3104
rect 8422 -3156 8434 -3104
rect 8486 -3156 8498 -3104
rect 8550 -3156 8562 -3104
rect 8614 -3156 8626 -3104
rect 8678 -3156 8690 -3104
rect 8742 -3156 8754 -3104
rect 8806 -3156 8818 -3104
rect 8870 -3156 8882 -3104
rect 8934 -3156 8960 -3104
rect 7980 -3172 8960 -3156
rect 7980 -3180 8316 -3172
rect 8577 -3180 8960 -3172
rect 9040 -3112 9120 -3080
rect 9240 -3081 10240 -3080
rect 9239 -3093 10240 -3081
rect 9040 -3116 9123 -3112
rect 9040 -3168 9055 -3116
rect 9107 -3168 9123 -3116
rect 9239 -3145 9264 -3093
rect 9316 -3145 9328 -3093
rect 9380 -3145 9392 -3093
rect 9444 -3145 9456 -3093
rect 9508 -3145 9520 -3093
rect 9572 -3145 9584 -3093
rect 9636 -3145 9648 -3093
rect 9700 -3145 9712 -3093
rect 9764 -3145 9776 -3093
rect 9828 -3145 9840 -3093
rect 9892 -3145 9904 -3093
rect 9956 -3145 9968 -3093
rect 10020 -3145 10032 -3093
rect 10084 -3145 10096 -3093
rect 10148 -3145 10160 -3093
rect 10212 -3145 10241 -3093
rect 9239 -3151 10241 -3145
rect 10300 -3104 10380 -3060
rect 11540 -2800 11640 -2680
rect 11758 -2621 12761 -2603
rect 11758 -2673 11789 -2621
rect 11841 -2673 11853 -2621
rect 11905 -2673 11917 -2621
rect 11969 -2673 11981 -2621
rect 12033 -2673 12045 -2621
rect 12097 -2673 12109 -2621
rect 12161 -2673 12173 -2621
rect 12225 -2673 12237 -2621
rect 12289 -2673 12301 -2621
rect 12353 -2673 12365 -2621
rect 12417 -2673 12429 -2621
rect 12481 -2673 12493 -2621
rect 12545 -2673 12557 -2621
rect 12609 -2673 12621 -2621
rect 12673 -2673 12685 -2621
rect 12737 -2673 12761 -2621
rect 11758 -2681 12761 -2673
rect 12840 -2680 12920 -2400
rect 13040 -2480 13540 -2400
rect 13660 -2434 13740 -2400
rect 13460 -2600 13520 -2480
rect 13040 -2680 13520 -2600
rect 12820 -2800 12920 -2680
rect 11540 -2822 11650 -2800
rect 11540 -2874 11574 -2822
rect 11626 -2874 11650 -2822
rect 11540 -2886 11650 -2874
rect 11540 -2938 11574 -2886
rect 11626 -2938 11650 -2886
rect 11540 -2960 11650 -2938
rect 12810 -2822 12920 -2800
rect 12810 -2874 12834 -2822
rect 12886 -2874 12920 -2822
rect 12810 -2886 12920 -2874
rect 12810 -2938 12834 -2886
rect 12886 -2938 12920 -2886
rect 12810 -2960 12920 -2938
rect 11540 -3080 11640 -2960
rect 12820 -3080 12920 -2960
rect 13420 -3080 13520 -2680
rect 13660 -2486 13672 -2434
rect 13724 -2486 13740 -2434
rect 9239 -3160 10240 -3151
rect 9040 -3172 9123 -3168
rect 9040 -3213 9120 -3172
rect 9240 -3180 10240 -3160
rect 10300 -3156 10313 -3104
rect 10365 -3156 10380 -3104
rect 10300 -3168 10380 -3156
rect 10300 -3220 10313 -3168
rect 10365 -3220 10380 -3168
rect 10500 -3108 11500 -3080
rect 10500 -3160 10553 -3108
rect 10605 -3160 10617 -3108
rect 10669 -3160 10681 -3108
rect 10733 -3160 10745 -3108
rect 10797 -3160 10809 -3108
rect 10861 -3160 10873 -3108
rect 10925 -3160 10937 -3108
rect 10989 -3160 11001 -3108
rect 11053 -3160 11065 -3108
rect 11117 -3160 11129 -3108
rect 11181 -3160 11193 -3108
rect 11245 -3160 11257 -3108
rect 11309 -3160 11321 -3108
rect 11373 -3160 11385 -3108
rect 11437 -3160 11500 -3108
rect 10500 -3180 11500 -3160
rect 10300 -3248 10380 -3220
rect 11560 -3221 11640 -3080
rect 11760 -3103 12760 -3080
rect 11760 -3155 11812 -3103
rect 11864 -3155 11876 -3103
rect 11928 -3155 11940 -3103
rect 11992 -3155 12004 -3103
rect 12056 -3155 12068 -3103
rect 12120 -3155 12132 -3103
rect 12184 -3155 12196 -3103
rect 12248 -3155 12260 -3103
rect 12312 -3155 12324 -3103
rect 12376 -3155 12388 -3103
rect 12440 -3155 12452 -3103
rect 12504 -3155 12516 -3103
rect 12568 -3155 12580 -3103
rect 12632 -3155 12644 -3103
rect 12696 -3155 12760 -3103
rect 11760 -3180 12760 -3155
rect 12840 -3240 12920 -3080
rect 13040 -3160 13520 -3080
rect 2280 -3360 2780 -3300
rect 2920 -3360 4080 -3300
rect 4200 -3360 5320 -3300
rect 5460 -3360 6580 -3280
rect 13460 -3300 13520 -3160
rect 6720 -3360 7920 -3300
rect 7960 -3360 9080 -3300
rect 9220 -3360 10360 -3300
rect 10480 -3360 11600 -3300
rect 11760 -3360 12860 -3300
rect 13020 -3360 13520 -3300
rect 2700 -3760 2780 -3360
rect 3960 -3760 4080 -3360
rect 5220 -3760 5320 -3360
rect 6480 -3760 6580 -3360
rect 7740 -3445 7920 -3360
rect 7740 -3479 7868 -3445
rect 7902 -3479 7920 -3445
rect 7740 -3517 7920 -3479
rect 7740 -3551 7868 -3517
rect 7902 -3551 7920 -3517
rect 7740 -3589 7920 -3551
rect 7740 -3623 7868 -3589
rect 7902 -3623 7920 -3589
rect 7740 -3661 7920 -3623
rect 7740 -3695 7868 -3661
rect 7902 -3695 7920 -3661
rect 7740 -3760 7920 -3695
rect 8980 -3760 9080 -3360
rect 10240 -3760 10360 -3360
rect 11480 -3760 11600 -3360
rect 12760 -3760 12860 -3360
rect 13420 -3760 13520 -3360
rect 2260 -3820 13520 -3760
rect 13550 -3112 13630 -3080
rect 13550 -3164 13564 -3112
rect 13616 -3164 13630 -3112
rect 5460 -3840 6580 -3820
rect 7740 -3840 7840 -3820
rect 2150 -4265 2163 -4213
rect 2215 -4265 2230 -4213
rect 2150 -4280 2230 -4265
rect 2260 -3892 2500 -3850
rect 2260 -3897 2419 -3892
rect 2260 -3949 2294 -3897
rect 2346 -3944 2419 -3897
rect 2471 -3944 2500 -3892
rect 2346 -3949 2500 -3944
rect 2260 -3956 2500 -3949
rect 2260 -3961 2419 -3956
rect 2260 -4013 2294 -3961
rect 2346 -4008 2419 -3961
rect 2471 -4008 2500 -3956
rect 2346 -4013 2500 -4008
rect 2020 -4598 2034 -4546
rect 2086 -4598 2100 -4546
rect 2020 -4610 2100 -4598
rect 2260 -4680 2500 -4013
rect 2100 -4740 2500 -4680
rect 2760 -3866 2840 -3850
rect 2760 -3918 2776 -3866
rect 2828 -3918 2840 -3866
rect 2760 -3930 2840 -3918
rect 2760 -3982 2776 -3930
rect 2828 -3982 2840 -3930
rect 2760 -3994 2840 -3982
rect 2760 -4046 2776 -3994
rect 2828 -4046 2840 -3994
rect 1890 -4772 2070 -4740
rect 1890 -4824 1914 -4772
rect 1966 -4824 2070 -4772
rect 1890 -4836 2070 -4824
rect 1890 -4888 1914 -4836
rect 1966 -4888 2070 -4836
rect 1890 -4940 2070 -4888
rect 2100 -4954 2500 -4950
rect 2100 -5006 2149 -4954
rect 2201 -5006 2289 -4954
rect 2341 -5006 2419 -4954
rect 2471 -5006 2500 -4954
rect 2100 -5010 2500 -5006
rect 2020 -5076 2730 -5060
rect 2020 -5078 2497 -5076
rect 2020 -5112 2048 -5078
rect 2082 -5112 2120 -5078
rect 2154 -5112 2192 -5078
rect 2226 -5112 2264 -5078
rect 2298 -5112 2336 -5078
rect 2370 -5112 2408 -5078
rect 2442 -5110 2497 -5078
rect 2531 -5110 2730 -5076
rect 2442 -5112 2730 -5110
rect 2020 -5160 2730 -5112
rect 2670 -6730 2730 -5160
rect 2760 -6234 2840 -4046
rect 9370 -3904 9450 -3850
rect 9370 -3956 9384 -3904
rect 9436 -3956 9450 -3904
rect 9370 -3994 9450 -3956
rect 9370 -4046 9384 -3994
rect 9436 -4046 9450 -3994
rect 2760 -6286 2774 -6234
rect 2826 -6286 2840 -6234
rect 2760 -6310 2840 -6286
rect 2870 -4104 2940 -4090
rect 2870 -4156 2879 -4104
rect 2931 -4156 2940 -4104
rect 2870 -4610 2940 -4156
rect 2670 -6746 2750 -6730
rect 2670 -6798 2681 -6746
rect 2733 -6798 2750 -6746
rect 2670 -6810 2750 -6798
rect 2670 -7410 2730 -6810
rect 2870 -6924 2950 -4610
rect 2870 -6976 2884 -6924
rect 2936 -6976 2950 -6924
rect 2870 -6990 2950 -6976
rect 2980 -4655 3060 -4640
rect 2980 -4707 2995 -4655
rect 3047 -4707 3060 -4655
rect 2980 -5526 3060 -4707
rect 3110 -4950 9230 -4870
rect 3510 -5350 3610 -4950
rect 4770 -5350 4850 -4950
rect 6010 -5350 6090 -4950
rect 7270 -5350 7350 -4950
rect 8510 -5350 8610 -4950
rect 9150 -5350 9230 -4950
rect 3110 -5410 3610 -5350
rect 3770 -5410 4850 -5350
rect 5010 -5410 6090 -5350
rect 6250 -5410 7350 -5350
rect 7490 -5410 8610 -5350
rect 8750 -5410 9230 -5350
rect 3510 -5510 3610 -5410
rect 2980 -5578 2996 -5526
rect 3048 -5578 3060 -5526
rect 2670 -7424 2770 -7410
rect 2670 -7476 2689 -7424
rect 2741 -7476 2770 -7424
rect 2670 -7490 2770 -7476
rect 2670 -8720 2730 -7490
rect 2980 -7604 3060 -5578
rect 3110 -5630 3610 -5510
rect 4030 -5547 4510 -5510
rect 4030 -5599 4126 -5547
rect 4178 -5599 4190 -5547
rect 4242 -5599 4254 -5547
rect 4306 -5599 4318 -5547
rect 4370 -5599 4382 -5547
rect 4434 -5599 4510 -5547
rect 4030 -5630 4510 -5599
rect 4790 -5516 4870 -5510
rect 4790 -5522 4873 -5516
rect 4790 -5574 4807 -5522
rect 4859 -5574 4873 -5522
rect 4790 -5579 4873 -5574
rect 5330 -5543 5810 -5510
rect 6050 -5516 6130 -5510
rect 3510 -6030 3610 -5630
rect 4790 -6030 4870 -5579
rect 5330 -5595 5413 -5543
rect 5465 -5595 5477 -5543
rect 5529 -5595 5541 -5543
rect 5593 -5595 5605 -5543
rect 5657 -5595 5669 -5543
rect 5721 -5595 5810 -5543
rect 6046 -5522 6130 -5516
rect 6046 -5574 6059 -5522
rect 6111 -5574 6130 -5522
rect 6046 -5579 6130 -5574
rect 5330 -5630 5810 -5595
rect 6050 -6030 6130 -5579
rect 6590 -5545 7070 -5510
rect 7290 -5515 7370 -5510
rect 6590 -5597 6693 -5545
rect 6745 -5597 6757 -5545
rect 6809 -5597 6821 -5545
rect 6873 -5597 6885 -5545
rect 6937 -5597 6949 -5545
rect 7001 -5597 7070 -5545
rect 7289 -5521 7370 -5515
rect 7289 -5573 7302 -5521
rect 7354 -5573 7370 -5521
rect 7289 -5578 7370 -5573
rect 6590 -5630 7070 -5597
rect 7290 -6030 7370 -5578
rect 7830 -5547 8310 -5510
rect 7830 -5599 7928 -5547
rect 7980 -5599 7992 -5547
rect 8044 -5599 8056 -5547
rect 8108 -5599 8120 -5547
rect 8172 -5599 8184 -5547
rect 8236 -5599 8310 -5547
rect 7830 -5630 8310 -5599
rect 8530 -5522 8610 -5510
rect 8530 -5574 8543 -5522
rect 8595 -5574 8610 -5522
rect 9150 -5570 9230 -5410
rect 3110 -6090 3610 -6030
rect 3510 -6250 3610 -6090
rect 3751 -6059 4757 -6035
rect 3751 -6111 3802 -6059
rect 3854 -6111 3866 -6059
rect 3918 -6111 3930 -6059
rect 3982 -6111 3994 -6059
rect 4046 -6111 4058 -6059
rect 4110 -6111 4122 -6059
rect 4174 -6111 4186 -6059
rect 4238 -6111 4250 -6059
rect 4302 -6111 4314 -6059
rect 4366 -6111 4378 -6059
rect 4430 -6111 4442 -6059
rect 4494 -6111 4506 -6059
rect 4558 -6111 4570 -6059
rect 4622 -6111 4634 -6059
rect 4686 -6111 4757 -6059
rect 3751 -6126 4757 -6111
rect 5005 -6063 6005 -6034
rect 5005 -6115 5031 -6063
rect 5083 -6115 5095 -6063
rect 5147 -6115 5159 -6063
rect 5211 -6115 5223 -6063
rect 5275 -6115 5287 -6063
rect 5339 -6115 5351 -6063
rect 5403 -6115 5415 -6063
rect 5467 -6115 5479 -6063
rect 5531 -6115 5543 -6063
rect 5595 -6115 5607 -6063
rect 5659 -6115 5671 -6063
rect 5723 -6115 5735 -6063
rect 5787 -6115 5799 -6063
rect 5851 -6115 5863 -6063
rect 5915 -6115 5927 -6063
rect 5979 -6115 6005 -6063
rect 5005 -6133 6005 -6115
rect 6249 -6061 7248 -6039
rect 6249 -6113 6275 -6061
rect 6327 -6113 6339 -6061
rect 6391 -6113 6403 -6061
rect 6455 -6113 6467 -6061
rect 6519 -6113 6531 -6061
rect 6583 -6113 6595 -6061
rect 6647 -6113 6659 -6061
rect 6711 -6113 6723 -6061
rect 6775 -6113 6787 -6061
rect 6839 -6113 6851 -6061
rect 6903 -6113 6915 -6061
rect 6967 -6113 6979 -6061
rect 7031 -6113 7043 -6061
rect 7095 -6113 7107 -6061
rect 7159 -6113 7171 -6061
rect 7223 -6113 7248 -6061
rect 6249 -6128 7248 -6113
rect 7490 -6066 8501 -6049
rect 7490 -6118 7513 -6066
rect 7565 -6118 7577 -6066
rect 7629 -6118 7641 -6066
rect 7693 -6118 7705 -6066
rect 7757 -6118 7769 -6066
rect 7821 -6118 7833 -6066
rect 7885 -6118 7897 -6066
rect 7949 -6118 7961 -6066
rect 8013 -6118 8025 -6066
rect 8077 -6118 8089 -6066
rect 8141 -6118 8153 -6066
rect 8205 -6118 8217 -6066
rect 8269 -6118 8281 -6066
rect 8333 -6118 8345 -6066
rect 8397 -6118 8409 -6066
rect 8461 -6118 8501 -6066
rect 7490 -6128 8501 -6118
rect 5090 -6227 5910 -6190
rect 3110 -6330 3610 -6250
rect 3761 -6250 4453 -6244
rect 3761 -6302 3793 -6250
rect 3845 -6302 3857 -6250
rect 3909 -6302 3921 -6250
rect 3973 -6302 3985 -6250
rect 4037 -6302 4049 -6250
rect 4101 -6302 4113 -6250
rect 4165 -6302 4177 -6250
rect 4229 -6302 4241 -6250
rect 4293 -6302 4305 -6250
rect 4357 -6302 4369 -6250
rect 4421 -6302 4453 -6250
rect 3761 -6307 4453 -6302
rect 5090 -6279 5124 -6227
rect 5176 -6279 5188 -6227
rect 5240 -6279 5252 -6227
rect 5304 -6279 5316 -6227
rect 5368 -6279 5380 -6227
rect 5432 -6279 5444 -6227
rect 5496 -6279 5508 -6227
rect 5560 -6279 5572 -6227
rect 5624 -6279 5636 -6227
rect 5688 -6279 5700 -6227
rect 5752 -6279 5764 -6227
rect 5816 -6279 5828 -6227
rect 5880 -6279 5910 -6227
rect 5090 -6310 5910 -6279
rect 6270 -6270 7450 -6210
rect 6270 -6310 7250 -6270
rect 7350 -6310 7450 -6270
rect 7672 -6233 8364 -6227
rect 7672 -6285 7704 -6233
rect 7756 -6285 7768 -6233
rect 7820 -6285 7832 -6233
rect 7884 -6285 7896 -6233
rect 7948 -6285 7960 -6233
rect 8012 -6285 8024 -6233
rect 8076 -6285 8088 -6233
rect 8140 -6285 8152 -6233
rect 8204 -6285 8216 -6233
rect 8268 -6285 8280 -6233
rect 8332 -6285 8364 -6233
rect 7672 -6290 8364 -6285
rect 3510 -6690 3610 -6330
rect 3110 -6770 3610 -6690
rect 4790 -6438 4870 -6310
rect 6050 -6312 6130 -6310
rect 6050 -6370 6197 -6312
rect 6050 -6422 6113 -6370
rect 6165 -6422 6197 -6370
rect 6050 -6434 6197 -6422
rect 4790 -6468 4879 -6438
rect 4790 -6520 4808 -6468
rect 4860 -6520 4879 -6468
rect 4790 -6532 4879 -6520
rect 4790 -6584 4808 -6532
rect 4860 -6584 4879 -6532
rect 4790 -6613 4879 -6584
rect 6050 -6486 6113 -6434
rect 6165 -6486 6197 -6434
rect 6050 -6498 6197 -6486
rect 6050 -6550 6113 -6498
rect 6165 -6550 6197 -6498
rect 6050 -6562 6197 -6550
rect 4790 -6710 4870 -6613
rect 6050 -6614 6113 -6562
rect 6165 -6614 6197 -6562
rect 6050 -6626 6197 -6614
rect 6050 -6678 6113 -6626
rect 6165 -6678 6197 -6626
rect 6050 -6710 6197 -6678
rect 7290 -6365 7450 -6310
rect 7290 -6417 7371 -6365
rect 7423 -6370 7450 -6365
rect 7423 -6417 7444 -6370
rect 7290 -6429 7444 -6417
rect 7290 -6481 7371 -6429
rect 7423 -6481 7444 -6429
rect 7290 -6493 7444 -6481
rect 7290 -6545 7371 -6493
rect 7423 -6545 7444 -6493
rect 7290 -6557 7444 -6545
rect 7290 -6609 7371 -6557
rect 7423 -6609 7444 -6557
rect 7290 -6621 7444 -6609
rect 7290 -6673 7371 -6621
rect 7423 -6673 7444 -6621
rect 7290 -6710 7444 -6673
rect 8530 -6710 8610 -5574
rect 8750 -5630 9250 -5570
rect 9150 -6030 9250 -5630
rect 8770 -6090 9250 -6030
rect 9150 -6250 9230 -6090
rect 8750 -6310 9230 -6250
rect 9150 -6710 9230 -6310
rect 3510 -6930 3610 -6770
rect 3751 -6742 4757 -6715
rect 3751 -6794 3781 -6742
rect 3833 -6794 3845 -6742
rect 3897 -6794 3909 -6742
rect 3961 -6794 3973 -6742
rect 4025 -6794 4037 -6742
rect 4089 -6794 4101 -6742
rect 4153 -6794 4165 -6742
rect 4217 -6794 4229 -6742
rect 4281 -6794 4293 -6742
rect 4345 -6794 4357 -6742
rect 4409 -6794 4421 -6742
rect 4473 -6794 4485 -6742
rect 4537 -6794 4549 -6742
rect 4601 -6794 4613 -6742
rect 4665 -6794 4677 -6742
rect 4729 -6794 4757 -6742
rect 3751 -6809 4757 -6794
rect 4990 -6748 5990 -6718
rect 4990 -6800 5024 -6748
rect 5076 -6800 5088 -6748
rect 5140 -6800 5152 -6748
rect 5204 -6800 5216 -6748
rect 5268 -6800 5280 -6748
rect 5332 -6800 5344 -6748
rect 5396 -6800 5408 -6748
rect 5460 -6800 5472 -6748
rect 5524 -6800 5536 -6748
rect 5588 -6800 5600 -6748
rect 5652 -6800 5664 -6748
rect 5716 -6800 5728 -6748
rect 5780 -6800 5792 -6748
rect 5844 -6800 5856 -6748
rect 5908 -6800 5920 -6748
rect 5972 -6800 5990 -6748
rect 4990 -6807 5990 -6800
rect 6050 -6890 6130 -6710
rect 6254 -6745 7251 -6711
rect 6254 -6797 6281 -6745
rect 6333 -6797 6345 -6745
rect 6397 -6797 6409 -6745
rect 6461 -6797 6473 -6745
rect 6525 -6797 6537 -6745
rect 6589 -6797 6601 -6745
rect 6653 -6797 6665 -6745
rect 6717 -6797 6729 -6745
rect 6781 -6797 6793 -6745
rect 6845 -6797 6857 -6745
rect 6909 -6797 6921 -6745
rect 6973 -6797 6985 -6745
rect 7037 -6797 7049 -6745
rect 7101 -6797 7113 -6745
rect 7165 -6797 7177 -6745
rect 7229 -6797 7251 -6745
rect 6254 -6814 7251 -6797
rect 3110 -6990 3610 -6930
rect 3760 -6926 4452 -6920
rect 3760 -6978 3792 -6926
rect 3844 -6978 3856 -6926
rect 3908 -6978 3920 -6926
rect 3972 -6978 3984 -6926
rect 4036 -6978 4048 -6926
rect 4100 -6978 4112 -6926
rect 4164 -6978 4176 -6926
rect 4228 -6978 4240 -6926
rect 4292 -6978 4304 -6926
rect 4356 -6978 4368 -6926
rect 4420 -6978 4452 -6926
rect 3760 -6983 4452 -6978
rect 4990 -6950 6130 -6890
rect 4990 -6990 5990 -6950
rect 3510 -7390 3610 -6990
rect 3110 -7450 3610 -7390
rect 2980 -7656 2994 -7604
rect 3046 -7656 3060 -7604
rect 3510 -7610 3610 -7450
rect 3751 -7421 4754 -7405
rect 3751 -7473 3775 -7421
rect 3827 -7473 3839 -7421
rect 3891 -7473 3903 -7421
rect 3955 -7473 3967 -7421
rect 4019 -7473 4031 -7421
rect 4083 -7473 4095 -7421
rect 4147 -7473 4159 -7421
rect 4211 -7473 4223 -7421
rect 4275 -7473 4287 -7421
rect 4339 -7473 4351 -7421
rect 4403 -7473 4415 -7421
rect 4467 -7473 4479 -7421
rect 4531 -7473 4543 -7421
rect 4595 -7473 4607 -7421
rect 4659 -7473 4671 -7421
rect 4723 -7473 4754 -7421
rect 3751 -7491 4754 -7473
rect 2980 -7670 3060 -7656
rect 3110 -7670 3610 -7610
rect 3890 -7596 4590 -7590
rect 3890 -7648 4112 -7596
rect 4164 -7648 4176 -7596
rect 4228 -7648 4240 -7596
rect 4292 -7648 4304 -7596
rect 4356 -7648 4590 -7596
rect 3890 -7650 4590 -7648
rect 4790 -7604 4870 -6990
rect 6050 -7390 6130 -6950
rect 6370 -6911 7190 -6870
rect 6370 -6963 6404 -6911
rect 6456 -6963 6468 -6911
rect 6520 -6963 6532 -6911
rect 6584 -6963 6596 -6911
rect 6648 -6963 6660 -6911
rect 6712 -6963 6724 -6911
rect 6776 -6963 6788 -6911
rect 6840 -6963 6852 -6911
rect 6904 -6963 6916 -6911
rect 6968 -6963 6980 -6911
rect 7032 -6963 7044 -6911
rect 7096 -6963 7108 -6911
rect 7160 -6963 7190 -6911
rect 6370 -6990 7190 -6963
rect 7290 -7390 7370 -6710
rect 7490 -6742 8487 -6722
rect 7490 -6794 7513 -6742
rect 7565 -6794 7577 -6742
rect 7629 -6794 7641 -6742
rect 7693 -6794 7705 -6742
rect 7757 -6794 7769 -6742
rect 7821 -6794 7833 -6742
rect 7885 -6794 7897 -6742
rect 7949 -6794 7961 -6742
rect 8013 -6794 8025 -6742
rect 8077 -6794 8089 -6742
rect 8141 -6794 8153 -6742
rect 8205 -6794 8217 -6742
rect 8269 -6794 8281 -6742
rect 8333 -6794 8345 -6742
rect 8397 -6794 8409 -6742
rect 8461 -6794 8487 -6742
rect 8750 -6770 9230 -6710
rect 7490 -6811 8487 -6794
rect 7501 -6925 8491 -6913
rect 7501 -6977 7659 -6925
rect 7711 -6977 7723 -6925
rect 7775 -6977 7787 -6925
rect 7839 -6977 7851 -6925
rect 7903 -6977 7915 -6925
rect 7967 -6977 7979 -6925
rect 8031 -6977 8043 -6925
rect 8095 -6977 8107 -6925
rect 8159 -6977 8171 -6925
rect 8223 -6977 8235 -6925
rect 8287 -6977 8491 -6925
rect 9150 -6930 9230 -6770
rect 7501 -6981 8491 -6977
rect 7627 -6982 8319 -6981
rect 8750 -6990 9230 -6930
rect 9370 -6924 9450 -4046
rect 9480 -4104 9640 -4090
rect 9480 -4156 9494 -4104
rect 9546 -4156 9574 -4104
rect 9626 -4156 9640 -4104
rect 9480 -4170 9640 -4156
rect 9480 -6234 9560 -4170
rect 13550 -4214 13630 -3164
rect 13550 -4266 13566 -4214
rect 13618 -4266 13630 -4214
rect 13550 -4280 13630 -4266
rect 13660 -4328 13740 -2486
rect 13660 -4380 13674 -4328
rect 13726 -4380 13740 -4328
rect 13660 -4390 13740 -4380
rect 13770 -4432 13850 -1778
rect 13770 -4484 13782 -4432
rect 13834 -4484 13850 -4432
rect 13770 -4500 13850 -4484
rect 13880 -4546 13960 -1104
rect 13880 -4598 13894 -4546
rect 13946 -4598 13960 -4546
rect 13880 -4610 13960 -4598
rect 9480 -6286 9494 -6234
rect 9546 -6286 9560 -6234
rect 9480 -6310 9560 -6286
rect 9590 -6064 9670 -6050
rect 9590 -6116 9604 -6064
rect 9656 -6116 9670 -6064
rect 9370 -6976 9385 -6924
rect 9437 -6976 9450 -6924
rect 9370 -6990 9450 -6976
rect 8530 -7058 8710 -6990
rect 8530 -7110 8624 -7058
rect 8676 -7110 8710 -7058
rect 8530 -7122 8710 -7110
rect 8530 -7174 8624 -7122
rect 8676 -7174 8710 -7122
rect 8530 -7186 8710 -7174
rect 8530 -7238 8624 -7186
rect 8676 -7238 8710 -7186
rect 8530 -7250 8710 -7238
rect 8530 -7302 8624 -7250
rect 8676 -7302 8710 -7250
rect 8530 -7390 8710 -7302
rect 9150 -7390 9230 -6990
rect 4991 -7421 5994 -7410
rect 4991 -7473 5014 -7421
rect 5066 -7473 5078 -7421
rect 5130 -7473 5142 -7421
rect 5194 -7473 5206 -7421
rect 5258 -7473 5270 -7421
rect 5322 -7473 5334 -7421
rect 5386 -7473 5398 -7421
rect 5450 -7473 5462 -7421
rect 5514 -7473 5526 -7421
rect 5578 -7473 5590 -7421
rect 5642 -7473 5654 -7421
rect 5706 -7473 5718 -7421
rect 5770 -7473 5782 -7421
rect 5834 -7473 5846 -7421
rect 5898 -7473 5910 -7421
rect 5962 -7473 5994 -7421
rect 4991 -7488 5994 -7473
rect 6233 -7425 7239 -7408
rect 6233 -7477 6256 -7425
rect 6308 -7477 6320 -7425
rect 6372 -7477 6384 -7425
rect 6436 -7477 6448 -7425
rect 6500 -7477 6512 -7425
rect 6564 -7477 6576 -7425
rect 6628 -7477 6640 -7425
rect 6692 -7477 6704 -7425
rect 6756 -7477 6768 -7425
rect 6820 -7477 6832 -7425
rect 6884 -7477 6896 -7425
rect 6948 -7477 6960 -7425
rect 7012 -7477 7024 -7425
rect 7076 -7477 7088 -7425
rect 7140 -7477 7152 -7425
rect 7204 -7477 7239 -7425
rect 6233 -7497 7239 -7477
rect 7495 -7422 8496 -7399
rect 7495 -7474 7516 -7422
rect 7568 -7474 7580 -7422
rect 7632 -7474 7644 -7422
rect 7696 -7474 7708 -7422
rect 7760 -7474 7772 -7422
rect 7824 -7474 7836 -7422
rect 7888 -7474 7900 -7422
rect 7952 -7474 7964 -7422
rect 8016 -7474 8028 -7422
rect 8080 -7474 8092 -7422
rect 8144 -7474 8156 -7422
rect 8208 -7474 8220 -7422
rect 8272 -7474 8284 -7422
rect 8336 -7474 8348 -7422
rect 8400 -7474 8412 -7422
rect 8464 -7474 8496 -7422
rect 8750 -7450 9230 -7390
rect 7495 -7497 8496 -7474
rect 3510 -8070 3610 -7670
rect 4790 -7656 4802 -7604
rect 4854 -7656 4870 -7604
rect 5170 -7596 5870 -7590
rect 5170 -7648 5340 -7596
rect 5392 -7648 5404 -7596
rect 5456 -7648 5468 -7596
rect 5520 -7648 5532 -7596
rect 5584 -7648 5870 -7596
rect 5170 -7650 5870 -7648
rect 6030 -7605 6110 -7590
rect 4790 -8050 4870 -7656
rect 6030 -7657 6041 -7605
rect 6093 -7657 6110 -7605
rect 6430 -7601 7130 -7590
rect 6430 -7650 6637 -7601
rect 6634 -7653 6637 -7650
rect 6689 -7653 6701 -7601
rect 6753 -7653 6765 -7601
rect 6817 -7653 6829 -7601
rect 6881 -7650 7130 -7601
rect 7270 -7611 7350 -7590
rect 6881 -7653 6885 -7650
rect 6634 -7655 6885 -7653
rect 6030 -8050 6110 -7657
rect 7270 -7663 7281 -7611
rect 7333 -7663 7350 -7611
rect 7650 -7597 8350 -7590
rect 7650 -7649 7905 -7597
rect 7957 -7649 7969 -7597
rect 8021 -7649 8033 -7597
rect 8085 -7649 8097 -7597
rect 8149 -7649 8350 -7597
rect 7650 -7650 8350 -7649
rect 8530 -7605 8610 -7590
rect 7902 -7651 8153 -7650
rect 7270 -8070 7350 -7663
rect 8530 -7657 8545 -7605
rect 8597 -7657 8610 -7605
rect 9150 -7610 9230 -7450
rect 8530 -8070 8610 -7657
rect 8750 -7670 9230 -7610
rect 9150 -8070 9230 -7670
rect 3110 -8130 3610 -8070
rect 2850 -8290 3060 -8280
rect 3510 -8290 3610 -8130
rect 3751 -8104 4752 -8090
rect 3751 -8156 3778 -8104
rect 3830 -8156 3842 -8104
rect 3894 -8156 3906 -8104
rect 3958 -8156 3970 -8104
rect 4022 -8156 4034 -8104
rect 4086 -8156 4098 -8104
rect 4150 -8156 4162 -8104
rect 4214 -8156 4226 -8104
rect 4278 -8156 4290 -8104
rect 4342 -8156 4354 -8104
rect 4406 -8156 4418 -8104
rect 4470 -8156 4482 -8104
rect 4534 -8156 4546 -8104
rect 4598 -8156 4610 -8104
rect 4662 -8156 4674 -8104
rect 4726 -8156 4752 -8104
rect 3751 -8170 4752 -8156
rect 4995 -8104 5992 -8083
rect 4995 -8156 5020 -8104
rect 5072 -8156 5084 -8104
rect 5136 -8156 5148 -8104
rect 5200 -8156 5212 -8104
rect 5264 -8156 5276 -8104
rect 5328 -8156 5340 -8104
rect 5392 -8156 5404 -8104
rect 5456 -8156 5468 -8104
rect 5520 -8156 5532 -8104
rect 5584 -8156 5596 -8104
rect 5648 -8156 5660 -8104
rect 5712 -8156 5724 -8104
rect 5776 -8156 5788 -8104
rect 5840 -8156 5852 -8104
rect 5904 -8156 5916 -8104
rect 5968 -8156 5992 -8104
rect 4995 -8173 5992 -8156
rect 6228 -8098 7232 -8083
rect 6228 -8150 6259 -8098
rect 6311 -8150 6323 -8098
rect 6375 -8150 6387 -8098
rect 6439 -8150 6451 -8098
rect 6503 -8150 6515 -8098
rect 6567 -8150 6579 -8098
rect 6631 -8150 6643 -8098
rect 6695 -8150 6707 -8098
rect 6759 -8150 6771 -8098
rect 6823 -8150 6835 -8098
rect 6887 -8150 6899 -8098
rect 6951 -8150 6963 -8098
rect 7015 -8150 7027 -8098
rect 7079 -8150 7091 -8098
rect 7143 -8150 7155 -8098
rect 7207 -8150 7232 -8098
rect 6228 -8170 7232 -8150
rect 7486 -8103 8496 -8082
rect 7486 -8155 7521 -8103
rect 7573 -8155 7585 -8103
rect 7637 -8155 7649 -8103
rect 7701 -8155 7713 -8103
rect 7765 -8155 7777 -8103
rect 7829 -8155 7841 -8103
rect 7893 -8155 7905 -8103
rect 7957 -8155 7969 -8103
rect 8021 -8155 8033 -8103
rect 8085 -8155 8097 -8103
rect 8149 -8155 8161 -8103
rect 8213 -8155 8225 -8103
rect 8277 -8155 8289 -8103
rect 8341 -8155 8353 -8103
rect 8405 -8155 8417 -8103
rect 8469 -8155 8496 -8103
rect 8750 -8130 9230 -8070
rect 7486 -8165 8496 -8155
rect 2850 -8296 3610 -8290
rect 2850 -8330 2993 -8296
rect 3027 -8330 3610 -8296
rect 9150 -8310 9230 -8130
rect 9590 -8104 9670 -6116
rect 9590 -8156 9604 -8104
rect 9656 -8156 9670 -8104
rect 9590 -8170 9670 -8156
rect 2850 -8331 3610 -8330
rect 2850 -8365 2883 -8331
rect 2917 -8365 3610 -8331
rect 2850 -8368 3610 -8365
rect 2850 -8402 2993 -8368
rect 3027 -8370 3610 -8368
rect 3750 -8370 4850 -8310
rect 5010 -8370 6090 -8310
rect 6250 -8370 7330 -8310
rect 7490 -8370 8570 -8310
rect 8750 -8370 9230 -8310
rect 3027 -8402 3130 -8370
rect 2850 -8403 3130 -8402
rect 2850 -8437 2883 -8403
rect 2917 -8437 3130 -8403
rect 2850 -8440 3130 -8437
rect 2850 -8474 2993 -8440
rect 3027 -8474 3130 -8440
rect 2850 -8475 3130 -8474
rect 2850 -8509 2883 -8475
rect 2917 -8509 3130 -8475
rect 2850 -8512 3130 -8509
rect 2850 -8546 2993 -8512
rect 3027 -8546 3130 -8512
rect 2850 -8547 3130 -8546
rect 2850 -8581 2883 -8547
rect 2917 -8581 3130 -8547
rect 2850 -8584 3130 -8581
rect 2850 -8618 2993 -8584
rect 3027 -8618 3130 -8584
rect 2850 -8619 3130 -8618
rect 2850 -8653 2883 -8619
rect 2917 -8653 3130 -8619
rect 2850 -8656 3130 -8653
rect 2850 -8690 2993 -8656
rect 3027 -8690 3130 -8656
rect 2850 -8691 3130 -8690
rect 2850 -8720 2883 -8691
rect 2670 -8725 2883 -8720
rect 2917 -8725 3130 -8691
rect 2670 -8728 3130 -8725
rect 2670 -8762 2993 -8728
rect 3027 -8750 3130 -8728
rect 3510 -8750 3610 -8370
rect 4770 -8750 4850 -8370
rect 6010 -8750 6090 -8370
rect 7250 -8750 7330 -8370
rect 8490 -8750 8570 -8370
rect 9150 -8750 9230 -8370
rect 3027 -8762 9230 -8750
rect 2670 -8763 9230 -8762
rect 2670 -8797 2883 -8763
rect 2917 -8797 9230 -8763
rect 2670 -8800 9230 -8797
rect 2670 -8834 2993 -8800
rect 3027 -8830 9230 -8800
rect 3027 -8834 3060 -8830
rect 2670 -8835 3060 -8834
rect 2670 -8869 2883 -8835
rect 2917 -8869 3060 -8835
rect 2670 -8890 3060 -8869
rect 2670 -8920 3030 -8890
<< via1 >>
rect 1914 224 1966 276
rect 1793 -1779 1845 -1727
rect 1682 -2477 1734 -2425
rect 1794 -4375 1846 -4323
rect 1681 -4485 1733 -4433
rect 3628 229 3680 281
rect 3692 229 3744 281
rect 3756 229 3808 281
rect 3820 229 3872 281
rect 6240 219 6292 271
rect 7824 229 7876 281
rect 7888 229 7940 281
rect 7952 229 8004 281
rect 8016 229 8068 281
rect 10539 226 10591 278
rect 2043 -605 2095 -553
rect 2951 -605 3003 -553
rect 3015 -605 3067 -553
rect 3079 -605 3131 -553
rect 3143 -605 3195 -553
rect 3207 -605 3259 -553
rect 3271 -605 3323 -553
rect 3335 -605 3387 -553
rect 3399 -605 3451 -553
rect 3463 -605 3515 -553
rect 3527 -605 3579 -553
rect 3591 -605 3643 -553
rect 3655 -605 3707 -553
rect 3719 -605 3771 -553
rect 3783 -605 3835 -553
rect 3847 -605 3899 -553
rect 4210 -609 4262 -557
rect 4274 -609 4326 -557
rect 4338 -609 4390 -557
rect 4402 -609 4454 -557
rect 4466 -609 4518 -557
rect 4530 -609 4582 -557
rect 4594 -609 4646 -557
rect 4658 -609 4710 -557
rect 4722 -609 4774 -557
rect 4786 -609 4838 -557
rect 4850 -609 4902 -557
rect 4914 -609 4966 -557
rect 4978 -609 5030 -557
rect 5042 -609 5094 -557
rect 5106 -609 5158 -557
rect 5474 -607 5526 -555
rect 5538 -607 5590 -555
rect 5602 -607 5654 -555
rect 5666 -607 5718 -555
rect 5730 -607 5782 -555
rect 5794 -607 5846 -555
rect 5858 -607 5910 -555
rect 5922 -607 5974 -555
rect 5986 -607 6038 -555
rect 6050 -607 6102 -555
rect 6114 -607 6166 -555
rect 6178 -607 6230 -555
rect 6242 -607 6294 -555
rect 6306 -607 6358 -555
rect 6370 -607 6422 -555
rect 6738 -611 6790 -559
rect 6802 -611 6854 -559
rect 6866 -611 6918 -559
rect 6930 -611 6982 -559
rect 6994 -611 7046 -559
rect 7058 -611 7110 -559
rect 7122 -611 7174 -559
rect 7186 -611 7238 -559
rect 7250 -611 7302 -559
rect 7314 -611 7366 -559
rect 7378 -611 7430 -559
rect 7442 -611 7494 -559
rect 7506 -611 7558 -559
rect 7570 -611 7622 -559
rect 7634 -611 7686 -559
rect 7993 -609 8045 -557
rect 8057 -609 8109 -557
rect 8121 -609 8173 -557
rect 8185 -609 8237 -557
rect 8249 -609 8301 -557
rect 8313 -609 8365 -557
rect 8377 -609 8429 -557
rect 8441 -609 8493 -557
rect 8505 -609 8557 -557
rect 8569 -609 8621 -557
rect 8633 -609 8685 -557
rect 8697 -609 8749 -557
rect 8761 -609 8813 -557
rect 8825 -609 8877 -557
rect 8889 -609 8941 -557
rect 3994 -814 4046 -762
rect 3994 -878 4046 -826
rect 5254 -814 5306 -762
rect 5254 -878 5306 -826
rect 6564 -760 6616 -708
rect 9264 -609 9316 -557
rect 9328 -609 9380 -557
rect 9392 -609 9444 -557
rect 9456 -609 9508 -557
rect 9520 -609 9572 -557
rect 9584 -609 9636 -557
rect 9648 -609 9700 -557
rect 9712 -609 9764 -557
rect 9776 -609 9828 -557
rect 9840 -609 9892 -557
rect 9904 -609 9956 -557
rect 9968 -609 10020 -557
rect 10032 -609 10084 -557
rect 10096 -609 10148 -557
rect 10160 -609 10212 -557
rect 10527 -612 10579 -560
rect 10591 -612 10643 -560
rect 10655 -612 10707 -560
rect 10719 -612 10771 -560
rect 10783 -612 10835 -560
rect 10847 -612 10899 -560
rect 10911 -612 10963 -560
rect 10975 -612 11027 -560
rect 11039 -612 11091 -560
rect 11103 -612 11155 -560
rect 11167 -612 11219 -560
rect 11231 -612 11283 -560
rect 11295 -612 11347 -560
rect 11359 -612 11411 -560
rect 11423 -612 11475 -560
rect 6564 -824 6616 -772
rect 6564 -888 6616 -836
rect 7774 -814 7826 -762
rect 7774 -878 7826 -826
rect 9034 -814 9086 -762
rect 9034 -878 9086 -826
rect 6564 -952 6616 -900
rect 11790 -612 11842 -560
rect 11854 -612 11906 -560
rect 11918 -612 11970 -560
rect 11982 -612 12034 -560
rect 12046 -612 12098 -560
rect 12110 -612 12162 -560
rect 12174 -612 12226 -560
rect 12238 -612 12290 -560
rect 12302 -612 12354 -560
rect 12366 -612 12418 -560
rect 12430 -612 12482 -560
rect 12494 -612 12546 -560
rect 12558 -612 12610 -560
rect 12622 -612 12674 -560
rect 12686 -612 12738 -560
rect 10356 -776 10408 -724
rect 10356 -840 10408 -788
rect 10356 -904 10408 -852
rect 10356 -968 10408 -916
rect 2162 -1107 2214 -1055
rect 2044 -1283 2096 -1231
rect 2044 -1967 2096 -1915
rect 2045 -2668 2097 -2616
rect 2032 -3158 2084 -3106
rect 2993 -1100 3045 -1048
rect 3057 -1100 3109 -1048
rect 3121 -1100 3173 -1048
rect 3185 -1100 3237 -1048
rect 3249 -1100 3301 -1048
rect 3313 -1100 3365 -1048
rect 3377 -1100 3429 -1048
rect 3441 -1100 3493 -1048
rect 3505 -1100 3557 -1048
rect 3569 -1100 3621 -1048
rect 3633 -1100 3685 -1048
rect 3697 -1100 3749 -1048
rect 3761 -1100 3813 -1048
rect 3825 -1100 3877 -1048
rect 2951 -1288 3003 -1236
rect 3015 -1288 3067 -1236
rect 3079 -1288 3131 -1236
rect 3143 -1288 3195 -1236
rect 3207 -1288 3259 -1236
rect 3271 -1288 3323 -1236
rect 3335 -1288 3387 -1236
rect 3399 -1288 3451 -1236
rect 3463 -1288 3515 -1236
rect 3527 -1288 3579 -1236
rect 3591 -1288 3643 -1236
rect 3655 -1288 3707 -1236
rect 3719 -1288 3771 -1236
rect 3783 -1288 3835 -1236
rect 3847 -1288 3899 -1236
rect 4239 -1102 4291 -1050
rect 4303 -1102 4355 -1050
rect 4367 -1102 4419 -1050
rect 4431 -1102 4483 -1050
rect 4495 -1102 4547 -1050
rect 4559 -1102 4611 -1050
rect 4623 -1102 4675 -1050
rect 4687 -1102 4739 -1050
rect 4751 -1102 4803 -1050
rect 4815 -1102 4867 -1050
rect 4879 -1102 4931 -1050
rect 4943 -1102 4995 -1050
rect 5007 -1102 5059 -1050
rect 5071 -1102 5123 -1050
rect 5275 -1106 5327 -1054
rect 5481 -1090 5533 -1038
rect 5545 -1090 5597 -1038
rect 5609 -1090 5661 -1038
rect 5673 -1090 5725 -1038
rect 5737 -1090 5789 -1038
rect 5801 -1090 5853 -1038
rect 5865 -1090 5917 -1038
rect 5929 -1090 5981 -1038
rect 5993 -1090 6045 -1038
rect 6057 -1090 6109 -1038
rect 6121 -1090 6173 -1038
rect 6185 -1090 6237 -1038
rect 6249 -1090 6301 -1038
rect 6313 -1090 6365 -1038
rect 6377 -1090 6429 -1038
rect 4220 -1294 4272 -1242
rect 4284 -1294 4336 -1242
rect 4348 -1294 4400 -1242
rect 4412 -1294 4464 -1242
rect 4476 -1294 4528 -1242
rect 4540 -1294 4592 -1242
rect 4604 -1294 4656 -1242
rect 4668 -1294 4720 -1242
rect 4732 -1294 4784 -1242
rect 4796 -1294 4848 -1242
rect 4860 -1294 4912 -1242
rect 4924 -1294 4976 -1242
rect 4988 -1294 5040 -1242
rect 5052 -1294 5104 -1242
rect 5116 -1294 5168 -1242
rect 6746 -1098 6798 -1046
rect 6810 -1098 6862 -1046
rect 6874 -1098 6926 -1046
rect 6938 -1098 6990 -1046
rect 7002 -1098 7054 -1046
rect 7066 -1098 7118 -1046
rect 7130 -1098 7182 -1046
rect 7194 -1098 7246 -1046
rect 7258 -1098 7310 -1046
rect 7322 -1098 7374 -1046
rect 7386 -1098 7438 -1046
rect 7450 -1098 7502 -1046
rect 7514 -1098 7566 -1046
rect 7578 -1098 7630 -1046
rect 3994 -1514 4046 -1462
rect 3994 -1578 4046 -1526
rect 5498 -1289 5550 -1237
rect 5562 -1289 5614 -1237
rect 5626 -1289 5678 -1237
rect 5690 -1289 5742 -1237
rect 5754 -1289 5806 -1237
rect 5818 -1289 5870 -1237
rect 5882 -1289 5934 -1237
rect 5946 -1289 5998 -1237
rect 6010 -1289 6062 -1237
rect 6074 -1289 6126 -1237
rect 6138 -1289 6190 -1237
rect 6202 -1289 6254 -1237
rect 6266 -1289 6318 -1237
rect 6330 -1289 6382 -1237
rect 6737 -1289 6789 -1237
rect 6801 -1289 6853 -1237
rect 6865 -1289 6917 -1237
rect 6929 -1289 6981 -1237
rect 6993 -1289 7045 -1237
rect 7057 -1289 7109 -1237
rect 7121 -1289 7173 -1237
rect 7185 -1289 7237 -1237
rect 7249 -1289 7301 -1237
rect 7313 -1289 7365 -1237
rect 7377 -1289 7429 -1237
rect 7441 -1289 7493 -1237
rect 7505 -1289 7557 -1237
rect 7569 -1289 7621 -1237
rect 7633 -1289 7685 -1237
rect 8004 -1098 8056 -1046
rect 8068 -1098 8120 -1046
rect 8132 -1098 8184 -1046
rect 8196 -1098 8248 -1046
rect 8260 -1098 8312 -1046
rect 8324 -1098 8376 -1046
rect 8388 -1098 8440 -1046
rect 8452 -1098 8504 -1046
rect 8516 -1098 8568 -1046
rect 8580 -1098 8632 -1046
rect 8644 -1098 8696 -1046
rect 8708 -1098 8760 -1046
rect 8772 -1098 8824 -1046
rect 8836 -1098 8888 -1046
rect 9053 -1106 9105 -1054
rect 9267 -1086 9319 -1034
rect 9331 -1086 9383 -1034
rect 9395 -1086 9447 -1034
rect 9459 -1086 9511 -1034
rect 9523 -1086 9575 -1034
rect 9587 -1086 9639 -1034
rect 9651 -1086 9703 -1034
rect 9715 -1086 9767 -1034
rect 9779 -1086 9831 -1034
rect 9843 -1086 9895 -1034
rect 9907 -1086 9959 -1034
rect 9971 -1086 10023 -1034
rect 10035 -1086 10087 -1034
rect 10099 -1086 10151 -1034
rect 10163 -1086 10215 -1034
rect 11574 -814 11626 -762
rect 11574 -878 11626 -826
rect 12834 -814 12886 -762
rect 12834 -878 12886 -826
rect 5274 -1514 5326 -1462
rect 5274 -1578 5326 -1526
rect 2974 -1784 3026 -1732
rect 3038 -1784 3090 -1732
rect 3102 -1784 3154 -1732
rect 3166 -1784 3218 -1732
rect 3230 -1784 3282 -1732
rect 3294 -1784 3346 -1732
rect 3358 -1784 3410 -1732
rect 3422 -1784 3474 -1732
rect 3486 -1784 3538 -1732
rect 3550 -1784 3602 -1732
rect 3614 -1784 3666 -1732
rect 3678 -1784 3730 -1732
rect 3742 -1784 3794 -1732
rect 3806 -1784 3858 -1732
rect 2950 -1963 3002 -1911
rect 3014 -1963 3066 -1911
rect 3078 -1963 3130 -1911
rect 3142 -1963 3194 -1911
rect 3206 -1963 3258 -1911
rect 3270 -1963 3322 -1911
rect 3334 -1963 3386 -1911
rect 3398 -1963 3450 -1911
rect 3462 -1963 3514 -1911
rect 3526 -1963 3578 -1911
rect 3590 -1963 3642 -1911
rect 3654 -1963 3706 -1911
rect 3718 -1963 3770 -1911
rect 3782 -1963 3834 -1911
rect 3846 -1963 3898 -1911
rect 4243 -1779 4295 -1727
rect 4307 -1779 4359 -1727
rect 4371 -1779 4423 -1727
rect 4435 -1779 4487 -1727
rect 4499 -1779 4551 -1727
rect 4563 -1779 4615 -1727
rect 4627 -1779 4679 -1727
rect 4691 -1779 4743 -1727
rect 4755 -1779 4807 -1727
rect 4819 -1779 4871 -1727
rect 4883 -1779 4935 -1727
rect 4947 -1779 4999 -1727
rect 5011 -1779 5063 -1727
rect 5075 -1779 5127 -1727
rect 4216 -1973 4268 -1921
rect 4280 -1973 4332 -1921
rect 4344 -1973 4396 -1921
rect 4408 -1973 4460 -1921
rect 4472 -1973 4524 -1921
rect 4536 -1973 4588 -1921
rect 4600 -1973 4652 -1921
rect 4664 -1973 4716 -1921
rect 4728 -1973 4780 -1921
rect 4792 -1973 4844 -1921
rect 4856 -1973 4908 -1921
rect 4920 -1973 4972 -1921
rect 4984 -1973 5036 -1921
rect 5048 -1973 5100 -1921
rect 5112 -1973 5164 -1921
rect 8020 -1283 8072 -1231
rect 8084 -1283 8136 -1231
rect 8148 -1283 8200 -1231
rect 8212 -1283 8264 -1231
rect 8276 -1283 8328 -1231
rect 8340 -1283 8392 -1231
rect 8404 -1283 8456 -1231
rect 8468 -1283 8520 -1231
rect 8532 -1283 8584 -1231
rect 8596 -1283 8648 -1231
rect 8660 -1283 8712 -1231
rect 8724 -1283 8776 -1231
rect 8788 -1283 8840 -1231
rect 8852 -1283 8904 -1231
rect 10548 -1101 10600 -1049
rect 10612 -1101 10664 -1049
rect 10676 -1101 10728 -1049
rect 10740 -1101 10792 -1049
rect 10804 -1101 10856 -1049
rect 10868 -1101 10920 -1049
rect 10932 -1101 10984 -1049
rect 10996 -1101 11048 -1049
rect 11060 -1101 11112 -1049
rect 11124 -1101 11176 -1049
rect 11188 -1101 11240 -1049
rect 11252 -1101 11304 -1049
rect 11316 -1101 11368 -1049
rect 11380 -1101 11432 -1049
rect 9283 -1295 9335 -1243
rect 9347 -1295 9399 -1243
rect 9411 -1295 9463 -1243
rect 9475 -1295 9527 -1243
rect 9539 -1295 9591 -1243
rect 9603 -1295 9655 -1243
rect 9667 -1295 9719 -1243
rect 9731 -1295 9783 -1243
rect 9795 -1295 9847 -1243
rect 9859 -1295 9911 -1243
rect 9923 -1295 9975 -1243
rect 9987 -1295 10039 -1243
rect 10051 -1295 10103 -1243
rect 10115 -1295 10167 -1243
rect 9054 -1514 9106 -1462
rect 9054 -1578 9106 -1526
rect 10525 -1295 10577 -1243
rect 10589 -1295 10641 -1243
rect 10653 -1295 10705 -1243
rect 10717 -1295 10769 -1243
rect 10781 -1295 10833 -1243
rect 10845 -1295 10897 -1243
rect 10909 -1295 10961 -1243
rect 10973 -1295 11025 -1243
rect 11037 -1295 11089 -1243
rect 11101 -1295 11153 -1243
rect 11165 -1295 11217 -1243
rect 11229 -1295 11281 -1243
rect 11293 -1295 11345 -1243
rect 11357 -1295 11409 -1243
rect 11421 -1295 11473 -1243
rect 11814 -1108 11866 -1056
rect 11878 -1108 11930 -1056
rect 11942 -1108 11994 -1056
rect 12006 -1108 12058 -1056
rect 12070 -1108 12122 -1056
rect 12134 -1108 12186 -1056
rect 12198 -1108 12250 -1056
rect 12262 -1108 12314 -1056
rect 12326 -1108 12378 -1056
rect 12390 -1108 12442 -1056
rect 12454 -1108 12506 -1056
rect 12518 -1108 12570 -1056
rect 12582 -1108 12634 -1056
rect 12646 -1108 12698 -1056
rect 11783 -1289 11835 -1237
rect 11847 -1289 11899 -1237
rect 11911 -1289 11963 -1237
rect 11975 -1289 12027 -1237
rect 12039 -1289 12091 -1237
rect 12103 -1289 12155 -1237
rect 12167 -1289 12219 -1237
rect 12231 -1289 12283 -1237
rect 12295 -1289 12347 -1237
rect 12359 -1289 12411 -1237
rect 12423 -1289 12475 -1237
rect 12487 -1289 12539 -1237
rect 12551 -1289 12603 -1237
rect 12615 -1289 12667 -1237
rect 12679 -1289 12731 -1237
rect 11574 -1514 11626 -1462
rect 11574 -1578 11626 -1526
rect 12834 -1514 12886 -1462
rect 12834 -1578 12886 -1526
rect 6762 -1789 6814 -1737
rect 6826 -1789 6878 -1737
rect 6890 -1789 6942 -1737
rect 6954 -1789 7006 -1737
rect 7018 -1789 7070 -1737
rect 7082 -1789 7134 -1737
rect 7146 -1789 7198 -1737
rect 7210 -1789 7262 -1737
rect 7274 -1789 7326 -1737
rect 7338 -1789 7390 -1737
rect 7402 -1789 7454 -1737
rect 7466 -1789 7518 -1737
rect 7530 -1789 7582 -1737
rect 7594 -1789 7646 -1737
rect 5480 -1965 5532 -1913
rect 5544 -1965 5596 -1913
rect 5608 -1965 5660 -1913
rect 5672 -1965 5724 -1913
rect 5736 -1965 5788 -1913
rect 5800 -1965 5852 -1913
rect 5864 -1965 5916 -1913
rect 5928 -1965 5980 -1913
rect 5992 -1965 6044 -1913
rect 6056 -1965 6108 -1913
rect 6120 -1965 6172 -1913
rect 6184 -1965 6236 -1913
rect 6248 -1965 6300 -1913
rect 6312 -1965 6364 -1913
rect 6376 -1965 6428 -1913
rect 6739 -1974 6791 -1922
rect 6803 -1974 6855 -1922
rect 6867 -1974 6919 -1922
rect 6931 -1974 6983 -1922
rect 6995 -1974 7047 -1922
rect 7059 -1974 7111 -1922
rect 7123 -1974 7175 -1922
rect 7187 -1974 7239 -1922
rect 7251 -1974 7303 -1922
rect 7315 -1974 7367 -1922
rect 7379 -1974 7431 -1922
rect 7443 -1974 7495 -1922
rect 7507 -1974 7559 -1922
rect 7571 -1974 7623 -1922
rect 7635 -1974 7687 -1922
rect 8021 -1786 8073 -1734
rect 8085 -1786 8137 -1734
rect 8149 -1786 8201 -1734
rect 8213 -1786 8265 -1734
rect 8277 -1786 8329 -1734
rect 8341 -1786 8393 -1734
rect 8405 -1786 8457 -1734
rect 8469 -1786 8521 -1734
rect 8533 -1786 8585 -1734
rect 8597 -1786 8649 -1734
rect 8661 -1786 8713 -1734
rect 8725 -1786 8777 -1734
rect 8789 -1786 8841 -1734
rect 8853 -1786 8905 -1734
rect 8000 -1975 8052 -1923
rect 8064 -1975 8116 -1923
rect 8128 -1975 8180 -1923
rect 8192 -1975 8244 -1923
rect 8256 -1975 8308 -1923
rect 8320 -1975 8372 -1923
rect 8384 -1975 8436 -1923
rect 8448 -1975 8500 -1923
rect 8512 -1975 8564 -1923
rect 8576 -1975 8628 -1923
rect 8640 -1975 8692 -1923
rect 8704 -1975 8756 -1923
rect 8768 -1975 8820 -1923
rect 8832 -1975 8884 -1923
rect 8896 -1975 8948 -1923
rect 10566 -1779 10618 -1727
rect 10630 -1779 10682 -1727
rect 10694 -1779 10746 -1727
rect 10758 -1779 10810 -1727
rect 10822 -1779 10874 -1727
rect 10886 -1779 10938 -1727
rect 10950 -1779 11002 -1727
rect 11014 -1779 11066 -1727
rect 11078 -1779 11130 -1727
rect 11142 -1779 11194 -1727
rect 11206 -1779 11258 -1727
rect 11270 -1779 11322 -1727
rect 11334 -1779 11386 -1727
rect 11398 -1779 11450 -1727
rect 9259 -1972 9311 -1920
rect 9323 -1972 9375 -1920
rect 9387 -1972 9439 -1920
rect 9451 -1972 9503 -1920
rect 9515 -1972 9567 -1920
rect 9579 -1972 9631 -1920
rect 9643 -1972 9695 -1920
rect 9707 -1972 9759 -1920
rect 9771 -1972 9823 -1920
rect 9835 -1972 9887 -1920
rect 9899 -1972 9951 -1920
rect 9963 -1972 10015 -1920
rect 10027 -1972 10079 -1920
rect 10091 -1972 10143 -1920
rect 10155 -1972 10207 -1920
rect 10521 -1976 10573 -1924
rect 10585 -1976 10637 -1924
rect 10649 -1976 10701 -1924
rect 10713 -1976 10765 -1924
rect 10777 -1976 10829 -1924
rect 10841 -1976 10893 -1924
rect 10905 -1976 10957 -1924
rect 10969 -1976 11021 -1924
rect 11033 -1976 11085 -1924
rect 11097 -1976 11149 -1924
rect 11161 -1976 11213 -1924
rect 11225 -1976 11277 -1924
rect 11289 -1976 11341 -1924
rect 11353 -1976 11405 -1924
rect 11417 -1976 11469 -1924
rect 11812 -1784 11864 -1732
rect 11876 -1784 11928 -1732
rect 11940 -1784 11992 -1732
rect 12004 -1784 12056 -1732
rect 12068 -1784 12120 -1732
rect 12132 -1784 12184 -1732
rect 12196 -1784 12248 -1732
rect 12260 -1784 12312 -1732
rect 12324 -1784 12376 -1732
rect 12388 -1784 12440 -1732
rect 12452 -1784 12504 -1732
rect 12516 -1784 12568 -1732
rect 12580 -1784 12632 -1732
rect 12644 -1784 12696 -1732
rect 11780 -1973 11832 -1921
rect 11844 -1973 11896 -1921
rect 11908 -1973 11960 -1921
rect 11972 -1973 12024 -1921
rect 12036 -1973 12088 -1921
rect 12100 -1973 12152 -1921
rect 12164 -1973 12216 -1921
rect 12228 -1973 12280 -1921
rect 12292 -1973 12344 -1921
rect 12356 -1973 12408 -1921
rect 12420 -1973 12472 -1921
rect 12484 -1973 12536 -1921
rect 12548 -1973 12600 -1921
rect 12612 -1973 12664 -1921
rect 12676 -1973 12728 -1921
rect 13892 -1104 13944 -1052
rect 13782 -1778 13834 -1726
rect 3994 -2214 4046 -2162
rect 3994 -2278 4046 -2226
rect 5254 -2214 5306 -2162
rect 5254 -2278 5306 -2226
rect 9054 -2214 9106 -2162
rect 9054 -2278 9106 -2226
rect 11574 -2214 11626 -2162
rect 11574 -2278 11626 -2226
rect 12834 -2214 12886 -2162
rect 12834 -2278 12886 -2226
rect 2974 -2477 3026 -2425
rect 3038 -2477 3090 -2425
rect 3102 -2477 3154 -2425
rect 3166 -2477 3218 -2425
rect 3230 -2477 3282 -2425
rect 3294 -2477 3346 -2425
rect 3358 -2477 3410 -2425
rect 3422 -2477 3474 -2425
rect 3486 -2477 3538 -2425
rect 3550 -2477 3602 -2425
rect 3614 -2477 3666 -2425
rect 3678 -2477 3730 -2425
rect 3742 -2477 3794 -2425
rect 3806 -2477 3858 -2425
rect 2947 -2664 2999 -2612
rect 3011 -2664 3063 -2612
rect 3075 -2664 3127 -2612
rect 3139 -2664 3191 -2612
rect 3203 -2664 3255 -2612
rect 3267 -2664 3319 -2612
rect 3331 -2664 3383 -2612
rect 3395 -2664 3447 -2612
rect 3459 -2664 3511 -2612
rect 3523 -2664 3575 -2612
rect 3587 -2664 3639 -2612
rect 3651 -2664 3703 -2612
rect 3715 -2664 3767 -2612
rect 3779 -2664 3831 -2612
rect 3843 -2664 3895 -2612
rect 4250 -2472 4302 -2420
rect 4314 -2472 4366 -2420
rect 4378 -2472 4430 -2420
rect 4442 -2472 4494 -2420
rect 4506 -2472 4558 -2420
rect 4570 -2472 4622 -2420
rect 4634 -2472 4686 -2420
rect 4698 -2472 4750 -2420
rect 4762 -2472 4814 -2420
rect 4826 -2472 4878 -2420
rect 4890 -2472 4942 -2420
rect 4954 -2472 5006 -2420
rect 5018 -2472 5070 -2420
rect 5082 -2472 5134 -2420
rect 4213 -2672 4265 -2620
rect 4277 -2672 4329 -2620
rect 4341 -2672 4393 -2620
rect 4405 -2672 4457 -2620
rect 4469 -2672 4521 -2620
rect 4533 -2672 4585 -2620
rect 4597 -2672 4649 -2620
rect 4661 -2672 4713 -2620
rect 4725 -2672 4777 -2620
rect 4789 -2672 4841 -2620
rect 4853 -2672 4905 -2620
rect 4917 -2672 4969 -2620
rect 4981 -2672 5033 -2620
rect 5045 -2672 5097 -2620
rect 5109 -2672 5161 -2620
rect 6759 -2467 6811 -2415
rect 6823 -2467 6875 -2415
rect 6887 -2467 6939 -2415
rect 6951 -2467 7003 -2415
rect 7015 -2467 7067 -2415
rect 7079 -2467 7131 -2415
rect 7143 -2467 7195 -2415
rect 7207 -2467 7259 -2415
rect 7271 -2467 7323 -2415
rect 7335 -2467 7387 -2415
rect 7399 -2467 7451 -2415
rect 7463 -2467 7515 -2415
rect 7527 -2467 7579 -2415
rect 7591 -2467 7643 -2415
rect 5479 -2672 5531 -2620
rect 5543 -2672 5595 -2620
rect 5607 -2672 5659 -2620
rect 5671 -2672 5723 -2620
rect 5735 -2672 5787 -2620
rect 5799 -2672 5851 -2620
rect 5863 -2672 5915 -2620
rect 5927 -2672 5979 -2620
rect 5991 -2672 6043 -2620
rect 6055 -2672 6107 -2620
rect 6119 -2672 6171 -2620
rect 6183 -2672 6235 -2620
rect 6247 -2672 6299 -2620
rect 6311 -2672 6363 -2620
rect 6375 -2672 6427 -2620
rect 6736 -2672 6788 -2620
rect 6800 -2672 6852 -2620
rect 6864 -2672 6916 -2620
rect 6928 -2672 6980 -2620
rect 6992 -2672 7044 -2620
rect 7056 -2672 7108 -2620
rect 7120 -2672 7172 -2620
rect 7184 -2672 7236 -2620
rect 7248 -2672 7300 -2620
rect 7312 -2672 7364 -2620
rect 7376 -2672 7428 -2620
rect 7440 -2672 7492 -2620
rect 7504 -2672 7556 -2620
rect 7568 -2672 7620 -2620
rect 7632 -2672 7684 -2620
rect 8009 -2458 8061 -2406
rect 8073 -2458 8125 -2406
rect 8137 -2458 8189 -2406
rect 8201 -2458 8253 -2406
rect 8265 -2458 8317 -2406
rect 8329 -2458 8381 -2406
rect 8393 -2458 8445 -2406
rect 8457 -2458 8509 -2406
rect 8521 -2458 8573 -2406
rect 8585 -2458 8637 -2406
rect 8649 -2458 8701 -2406
rect 8713 -2458 8765 -2406
rect 8777 -2458 8829 -2406
rect 8841 -2458 8893 -2406
rect 3994 -2874 4046 -2822
rect 3994 -2938 4046 -2886
rect 5254 -2874 5306 -2822
rect 5254 -2938 5306 -2886
rect 8004 -2672 8056 -2620
rect 8068 -2672 8120 -2620
rect 8132 -2672 8184 -2620
rect 8196 -2672 8248 -2620
rect 8260 -2672 8312 -2620
rect 8324 -2672 8376 -2620
rect 8388 -2672 8440 -2620
rect 8452 -2672 8504 -2620
rect 8516 -2672 8568 -2620
rect 8580 -2672 8632 -2620
rect 8644 -2672 8696 -2620
rect 8708 -2672 8760 -2620
rect 8772 -2672 8824 -2620
rect 8836 -2672 8888 -2620
rect 8900 -2672 8952 -2620
rect 9264 -2669 9316 -2617
rect 9328 -2669 9380 -2617
rect 9392 -2669 9444 -2617
rect 9456 -2669 9508 -2617
rect 9520 -2669 9572 -2617
rect 9584 -2669 9636 -2617
rect 9648 -2669 9700 -2617
rect 9712 -2669 9764 -2617
rect 9776 -2669 9828 -2617
rect 9840 -2669 9892 -2617
rect 9904 -2669 9956 -2617
rect 9968 -2669 10020 -2617
rect 10032 -2669 10084 -2617
rect 10096 -2669 10148 -2617
rect 10160 -2669 10212 -2617
rect 10564 -2476 10616 -2424
rect 10628 -2476 10680 -2424
rect 10692 -2476 10744 -2424
rect 10756 -2476 10808 -2424
rect 10820 -2476 10872 -2424
rect 10884 -2476 10936 -2424
rect 10948 -2476 11000 -2424
rect 11012 -2476 11064 -2424
rect 11076 -2476 11128 -2424
rect 11140 -2476 11192 -2424
rect 11204 -2476 11256 -2424
rect 11268 -2476 11320 -2424
rect 11332 -2476 11384 -2424
rect 11396 -2476 11448 -2424
rect 9054 -2874 9106 -2822
rect 9054 -2938 9106 -2886
rect 10525 -2668 10577 -2616
rect 10589 -2668 10641 -2616
rect 10653 -2668 10705 -2616
rect 10717 -2668 10769 -2616
rect 10781 -2668 10833 -2616
rect 10845 -2668 10897 -2616
rect 10909 -2668 10961 -2616
rect 10973 -2668 11025 -2616
rect 11037 -2668 11089 -2616
rect 11101 -2668 11153 -2616
rect 11165 -2668 11217 -2616
rect 11229 -2668 11281 -2616
rect 11293 -2668 11345 -2616
rect 11357 -2668 11409 -2616
rect 11421 -2668 11473 -2616
rect 11812 -2481 11864 -2429
rect 11876 -2481 11928 -2429
rect 11940 -2481 11992 -2429
rect 12004 -2481 12056 -2429
rect 12068 -2481 12120 -2429
rect 12132 -2481 12184 -2429
rect 12196 -2481 12248 -2429
rect 12260 -2481 12312 -2429
rect 12324 -2481 12376 -2429
rect 12388 -2481 12440 -2429
rect 12452 -2481 12504 -2429
rect 12516 -2481 12568 -2429
rect 12580 -2481 12632 -2429
rect 12644 -2481 12696 -2429
rect 2969 -3160 3021 -3108
rect 3033 -3160 3085 -3108
rect 3097 -3160 3149 -3108
rect 3161 -3160 3213 -3108
rect 3225 -3160 3277 -3108
rect 3289 -3160 3341 -3108
rect 3353 -3160 3405 -3108
rect 3417 -3160 3469 -3108
rect 3481 -3160 3533 -3108
rect 3545 -3160 3597 -3108
rect 3609 -3160 3661 -3108
rect 3673 -3160 3725 -3108
rect 3737 -3160 3789 -3108
rect 3801 -3160 3853 -3108
rect 4248 -3167 4300 -3115
rect 4312 -3167 4364 -3115
rect 4376 -3167 4428 -3115
rect 4440 -3167 4492 -3115
rect 4504 -3167 4556 -3115
rect 4568 -3167 4620 -3115
rect 4632 -3167 4684 -3115
rect 4696 -3167 4748 -3115
rect 4760 -3167 4812 -3115
rect 4824 -3167 4876 -3115
rect 4888 -3167 4940 -3115
rect 4952 -3167 5004 -3115
rect 5016 -3167 5068 -3115
rect 5080 -3167 5132 -3115
rect 5273 -3169 5325 -3117
rect 5474 -3148 5526 -3096
rect 5538 -3148 5590 -3096
rect 5602 -3148 5654 -3096
rect 5666 -3148 5718 -3096
rect 5730 -3148 5782 -3096
rect 5794 -3148 5846 -3096
rect 5858 -3148 5910 -3096
rect 5922 -3148 5974 -3096
rect 5986 -3148 6038 -3096
rect 6050 -3148 6102 -3096
rect 6114 -3148 6166 -3096
rect 6178 -3148 6230 -3096
rect 6242 -3148 6294 -3096
rect 6306 -3148 6358 -3096
rect 6370 -3148 6422 -3096
rect 6726 -3156 6778 -3104
rect 6790 -3156 6842 -3104
rect 6854 -3156 6906 -3104
rect 6918 -3156 6970 -3104
rect 6982 -3156 7034 -3104
rect 7046 -3156 7098 -3104
rect 7110 -3156 7162 -3104
rect 7174 -3156 7226 -3104
rect 7238 -3156 7290 -3104
rect 7302 -3156 7354 -3104
rect 7366 -3156 7418 -3104
rect 7430 -3156 7482 -3104
rect 7494 -3156 7546 -3104
rect 7558 -3156 7610 -3104
rect 7622 -3156 7674 -3104
rect 7986 -3156 8038 -3104
rect 8050 -3156 8102 -3104
rect 8114 -3156 8166 -3104
rect 8178 -3156 8230 -3104
rect 8242 -3156 8294 -3104
rect 8306 -3156 8358 -3104
rect 8370 -3156 8422 -3104
rect 8434 -3156 8486 -3104
rect 8498 -3156 8550 -3104
rect 8562 -3156 8614 -3104
rect 8626 -3156 8678 -3104
rect 8690 -3156 8742 -3104
rect 8754 -3156 8806 -3104
rect 8818 -3156 8870 -3104
rect 8882 -3156 8934 -3104
rect 9055 -3168 9107 -3116
rect 9264 -3145 9316 -3093
rect 9328 -3145 9380 -3093
rect 9392 -3145 9444 -3093
rect 9456 -3145 9508 -3093
rect 9520 -3145 9572 -3093
rect 9584 -3145 9636 -3093
rect 9648 -3145 9700 -3093
rect 9712 -3145 9764 -3093
rect 9776 -3145 9828 -3093
rect 9840 -3145 9892 -3093
rect 9904 -3145 9956 -3093
rect 9968 -3145 10020 -3093
rect 10032 -3145 10084 -3093
rect 10096 -3145 10148 -3093
rect 10160 -3145 10212 -3093
rect 11789 -2673 11841 -2621
rect 11853 -2673 11905 -2621
rect 11917 -2673 11969 -2621
rect 11981 -2673 12033 -2621
rect 12045 -2673 12097 -2621
rect 12109 -2673 12161 -2621
rect 12173 -2673 12225 -2621
rect 12237 -2673 12289 -2621
rect 12301 -2673 12353 -2621
rect 12365 -2673 12417 -2621
rect 12429 -2673 12481 -2621
rect 12493 -2673 12545 -2621
rect 12557 -2673 12609 -2621
rect 12621 -2673 12673 -2621
rect 12685 -2673 12737 -2621
rect 11574 -2874 11626 -2822
rect 11574 -2938 11626 -2886
rect 12834 -2874 12886 -2822
rect 12834 -2938 12886 -2886
rect 13672 -2486 13724 -2434
rect 10313 -3156 10365 -3104
rect 10313 -3220 10365 -3168
rect 10553 -3160 10605 -3108
rect 10617 -3160 10669 -3108
rect 10681 -3160 10733 -3108
rect 10745 -3160 10797 -3108
rect 10809 -3160 10861 -3108
rect 10873 -3160 10925 -3108
rect 10937 -3160 10989 -3108
rect 11001 -3160 11053 -3108
rect 11065 -3160 11117 -3108
rect 11129 -3160 11181 -3108
rect 11193 -3160 11245 -3108
rect 11257 -3160 11309 -3108
rect 11321 -3160 11373 -3108
rect 11385 -3160 11437 -3108
rect 11812 -3155 11864 -3103
rect 11876 -3155 11928 -3103
rect 11940 -3155 11992 -3103
rect 12004 -3155 12056 -3103
rect 12068 -3155 12120 -3103
rect 12132 -3155 12184 -3103
rect 12196 -3155 12248 -3103
rect 12260 -3155 12312 -3103
rect 12324 -3155 12376 -3103
rect 12388 -3155 12440 -3103
rect 12452 -3155 12504 -3103
rect 12516 -3155 12568 -3103
rect 12580 -3155 12632 -3103
rect 12644 -3155 12696 -3103
rect 13564 -3164 13616 -3112
rect 2163 -4265 2215 -4213
rect 2294 -3949 2346 -3897
rect 2419 -3944 2471 -3892
rect 2294 -4013 2346 -3961
rect 2419 -4008 2471 -3956
rect 2034 -4598 2086 -4546
rect 2776 -3918 2828 -3866
rect 2776 -3982 2828 -3930
rect 2776 -4046 2828 -3994
rect 1914 -4824 1966 -4772
rect 1914 -4888 1966 -4836
rect 2149 -5006 2201 -4954
rect 2289 -5006 2341 -4954
rect 2419 -5006 2471 -4954
rect 9384 -3956 9436 -3904
rect 9384 -4046 9436 -3994
rect 2774 -6286 2826 -6234
rect 2879 -4156 2931 -4104
rect 2681 -6798 2733 -6746
rect 2884 -6976 2936 -6924
rect 2995 -4707 3047 -4655
rect 2996 -5578 3048 -5526
rect 2689 -7476 2741 -7424
rect 4126 -5599 4178 -5547
rect 4190 -5599 4242 -5547
rect 4254 -5599 4306 -5547
rect 4318 -5599 4370 -5547
rect 4382 -5599 4434 -5547
rect 4807 -5574 4859 -5522
rect 5413 -5595 5465 -5543
rect 5477 -5595 5529 -5543
rect 5541 -5595 5593 -5543
rect 5605 -5595 5657 -5543
rect 5669 -5595 5721 -5543
rect 6059 -5574 6111 -5522
rect 6693 -5597 6745 -5545
rect 6757 -5597 6809 -5545
rect 6821 -5597 6873 -5545
rect 6885 -5597 6937 -5545
rect 6949 -5597 7001 -5545
rect 7302 -5573 7354 -5521
rect 7928 -5599 7980 -5547
rect 7992 -5599 8044 -5547
rect 8056 -5599 8108 -5547
rect 8120 -5599 8172 -5547
rect 8184 -5599 8236 -5547
rect 8543 -5574 8595 -5522
rect 3802 -6111 3854 -6059
rect 3866 -6111 3918 -6059
rect 3930 -6111 3982 -6059
rect 3994 -6111 4046 -6059
rect 4058 -6111 4110 -6059
rect 4122 -6111 4174 -6059
rect 4186 -6111 4238 -6059
rect 4250 -6111 4302 -6059
rect 4314 -6111 4366 -6059
rect 4378 -6111 4430 -6059
rect 4442 -6111 4494 -6059
rect 4506 -6111 4558 -6059
rect 4570 -6111 4622 -6059
rect 4634 -6111 4686 -6059
rect 5031 -6115 5083 -6063
rect 5095 -6115 5147 -6063
rect 5159 -6115 5211 -6063
rect 5223 -6115 5275 -6063
rect 5287 -6115 5339 -6063
rect 5351 -6115 5403 -6063
rect 5415 -6115 5467 -6063
rect 5479 -6115 5531 -6063
rect 5543 -6115 5595 -6063
rect 5607 -6115 5659 -6063
rect 5671 -6115 5723 -6063
rect 5735 -6115 5787 -6063
rect 5799 -6115 5851 -6063
rect 5863 -6115 5915 -6063
rect 5927 -6115 5979 -6063
rect 6275 -6113 6327 -6061
rect 6339 -6113 6391 -6061
rect 6403 -6113 6455 -6061
rect 6467 -6113 6519 -6061
rect 6531 -6113 6583 -6061
rect 6595 -6113 6647 -6061
rect 6659 -6113 6711 -6061
rect 6723 -6113 6775 -6061
rect 6787 -6113 6839 -6061
rect 6851 -6113 6903 -6061
rect 6915 -6113 6967 -6061
rect 6979 -6113 7031 -6061
rect 7043 -6113 7095 -6061
rect 7107 -6113 7159 -6061
rect 7171 -6113 7223 -6061
rect 7513 -6118 7565 -6066
rect 7577 -6118 7629 -6066
rect 7641 -6118 7693 -6066
rect 7705 -6118 7757 -6066
rect 7769 -6118 7821 -6066
rect 7833 -6118 7885 -6066
rect 7897 -6118 7949 -6066
rect 7961 -6118 8013 -6066
rect 8025 -6118 8077 -6066
rect 8089 -6118 8141 -6066
rect 8153 -6118 8205 -6066
rect 8217 -6118 8269 -6066
rect 8281 -6118 8333 -6066
rect 8345 -6118 8397 -6066
rect 8409 -6118 8461 -6066
rect 3793 -6302 3845 -6250
rect 3857 -6302 3909 -6250
rect 3921 -6302 3973 -6250
rect 3985 -6302 4037 -6250
rect 4049 -6302 4101 -6250
rect 4113 -6302 4165 -6250
rect 4177 -6302 4229 -6250
rect 4241 -6302 4293 -6250
rect 4305 -6302 4357 -6250
rect 4369 -6302 4421 -6250
rect 5124 -6279 5176 -6227
rect 5188 -6279 5240 -6227
rect 5252 -6279 5304 -6227
rect 5316 -6279 5368 -6227
rect 5380 -6279 5432 -6227
rect 5444 -6279 5496 -6227
rect 5508 -6279 5560 -6227
rect 5572 -6279 5624 -6227
rect 5636 -6279 5688 -6227
rect 5700 -6279 5752 -6227
rect 5764 -6279 5816 -6227
rect 5828 -6279 5880 -6227
rect 7704 -6285 7756 -6233
rect 7768 -6285 7820 -6233
rect 7832 -6285 7884 -6233
rect 7896 -6285 7948 -6233
rect 7960 -6285 8012 -6233
rect 8024 -6285 8076 -6233
rect 8088 -6285 8140 -6233
rect 8152 -6285 8204 -6233
rect 8216 -6285 8268 -6233
rect 8280 -6285 8332 -6233
rect 6113 -6422 6165 -6370
rect 4808 -6520 4860 -6468
rect 4808 -6584 4860 -6532
rect 6113 -6486 6165 -6434
rect 6113 -6550 6165 -6498
rect 6113 -6614 6165 -6562
rect 6113 -6678 6165 -6626
rect 7371 -6417 7423 -6365
rect 7371 -6481 7423 -6429
rect 7371 -6545 7423 -6493
rect 7371 -6609 7423 -6557
rect 7371 -6673 7423 -6621
rect 3781 -6794 3833 -6742
rect 3845 -6794 3897 -6742
rect 3909 -6794 3961 -6742
rect 3973 -6794 4025 -6742
rect 4037 -6794 4089 -6742
rect 4101 -6794 4153 -6742
rect 4165 -6794 4217 -6742
rect 4229 -6794 4281 -6742
rect 4293 -6794 4345 -6742
rect 4357 -6794 4409 -6742
rect 4421 -6794 4473 -6742
rect 4485 -6794 4537 -6742
rect 4549 -6794 4601 -6742
rect 4613 -6794 4665 -6742
rect 4677 -6794 4729 -6742
rect 5024 -6800 5076 -6748
rect 5088 -6800 5140 -6748
rect 5152 -6800 5204 -6748
rect 5216 -6800 5268 -6748
rect 5280 -6800 5332 -6748
rect 5344 -6800 5396 -6748
rect 5408 -6800 5460 -6748
rect 5472 -6800 5524 -6748
rect 5536 -6800 5588 -6748
rect 5600 -6800 5652 -6748
rect 5664 -6800 5716 -6748
rect 5728 -6800 5780 -6748
rect 5792 -6800 5844 -6748
rect 5856 -6800 5908 -6748
rect 5920 -6800 5972 -6748
rect 6281 -6797 6333 -6745
rect 6345 -6797 6397 -6745
rect 6409 -6797 6461 -6745
rect 6473 -6797 6525 -6745
rect 6537 -6797 6589 -6745
rect 6601 -6797 6653 -6745
rect 6665 -6797 6717 -6745
rect 6729 -6797 6781 -6745
rect 6793 -6797 6845 -6745
rect 6857 -6797 6909 -6745
rect 6921 -6797 6973 -6745
rect 6985 -6797 7037 -6745
rect 7049 -6797 7101 -6745
rect 7113 -6797 7165 -6745
rect 7177 -6797 7229 -6745
rect 3792 -6978 3844 -6926
rect 3856 -6978 3908 -6926
rect 3920 -6978 3972 -6926
rect 3984 -6978 4036 -6926
rect 4048 -6978 4100 -6926
rect 4112 -6978 4164 -6926
rect 4176 -6978 4228 -6926
rect 4240 -6978 4292 -6926
rect 4304 -6978 4356 -6926
rect 4368 -6978 4420 -6926
rect 2994 -7656 3046 -7604
rect 3775 -7473 3827 -7421
rect 3839 -7473 3891 -7421
rect 3903 -7473 3955 -7421
rect 3967 -7473 4019 -7421
rect 4031 -7473 4083 -7421
rect 4095 -7473 4147 -7421
rect 4159 -7473 4211 -7421
rect 4223 -7473 4275 -7421
rect 4287 -7473 4339 -7421
rect 4351 -7473 4403 -7421
rect 4415 -7473 4467 -7421
rect 4479 -7473 4531 -7421
rect 4543 -7473 4595 -7421
rect 4607 -7473 4659 -7421
rect 4671 -7473 4723 -7421
rect 4112 -7648 4164 -7596
rect 4176 -7648 4228 -7596
rect 4240 -7648 4292 -7596
rect 4304 -7648 4356 -7596
rect 6404 -6963 6456 -6911
rect 6468 -6963 6520 -6911
rect 6532 -6963 6584 -6911
rect 6596 -6963 6648 -6911
rect 6660 -6963 6712 -6911
rect 6724 -6963 6776 -6911
rect 6788 -6963 6840 -6911
rect 6852 -6963 6904 -6911
rect 6916 -6963 6968 -6911
rect 6980 -6963 7032 -6911
rect 7044 -6963 7096 -6911
rect 7108 -6963 7160 -6911
rect 7513 -6794 7565 -6742
rect 7577 -6794 7629 -6742
rect 7641 -6794 7693 -6742
rect 7705 -6794 7757 -6742
rect 7769 -6794 7821 -6742
rect 7833 -6794 7885 -6742
rect 7897 -6794 7949 -6742
rect 7961 -6794 8013 -6742
rect 8025 -6794 8077 -6742
rect 8089 -6794 8141 -6742
rect 8153 -6794 8205 -6742
rect 8217 -6794 8269 -6742
rect 8281 -6794 8333 -6742
rect 8345 -6794 8397 -6742
rect 8409 -6794 8461 -6742
rect 7659 -6977 7711 -6925
rect 7723 -6977 7775 -6925
rect 7787 -6977 7839 -6925
rect 7851 -6977 7903 -6925
rect 7915 -6977 7967 -6925
rect 7979 -6977 8031 -6925
rect 8043 -6977 8095 -6925
rect 8107 -6977 8159 -6925
rect 8171 -6977 8223 -6925
rect 8235 -6977 8287 -6925
rect 9494 -4156 9546 -4104
rect 9574 -4156 9626 -4104
rect 13566 -4266 13618 -4214
rect 13674 -4380 13726 -4328
rect 13782 -4484 13834 -4432
rect 13894 -4598 13946 -4546
rect 9494 -6286 9546 -6234
rect 9604 -6116 9656 -6064
rect 9385 -6976 9437 -6924
rect 8624 -7110 8676 -7058
rect 8624 -7174 8676 -7122
rect 8624 -7238 8676 -7186
rect 8624 -7302 8676 -7250
rect 5014 -7473 5066 -7421
rect 5078 -7473 5130 -7421
rect 5142 -7473 5194 -7421
rect 5206 -7473 5258 -7421
rect 5270 -7473 5322 -7421
rect 5334 -7473 5386 -7421
rect 5398 -7473 5450 -7421
rect 5462 -7473 5514 -7421
rect 5526 -7473 5578 -7421
rect 5590 -7473 5642 -7421
rect 5654 -7473 5706 -7421
rect 5718 -7473 5770 -7421
rect 5782 -7473 5834 -7421
rect 5846 -7473 5898 -7421
rect 5910 -7473 5962 -7421
rect 6256 -7477 6308 -7425
rect 6320 -7477 6372 -7425
rect 6384 -7477 6436 -7425
rect 6448 -7477 6500 -7425
rect 6512 -7477 6564 -7425
rect 6576 -7477 6628 -7425
rect 6640 -7477 6692 -7425
rect 6704 -7477 6756 -7425
rect 6768 -7477 6820 -7425
rect 6832 -7477 6884 -7425
rect 6896 -7477 6948 -7425
rect 6960 -7477 7012 -7425
rect 7024 -7477 7076 -7425
rect 7088 -7477 7140 -7425
rect 7152 -7477 7204 -7425
rect 7516 -7474 7568 -7422
rect 7580 -7474 7632 -7422
rect 7644 -7474 7696 -7422
rect 7708 -7474 7760 -7422
rect 7772 -7474 7824 -7422
rect 7836 -7474 7888 -7422
rect 7900 -7474 7952 -7422
rect 7964 -7474 8016 -7422
rect 8028 -7474 8080 -7422
rect 8092 -7474 8144 -7422
rect 8156 -7474 8208 -7422
rect 8220 -7474 8272 -7422
rect 8284 -7474 8336 -7422
rect 8348 -7474 8400 -7422
rect 8412 -7474 8464 -7422
rect 4802 -7656 4854 -7604
rect 5340 -7648 5392 -7596
rect 5404 -7648 5456 -7596
rect 5468 -7648 5520 -7596
rect 5532 -7648 5584 -7596
rect 6041 -7657 6093 -7605
rect 6637 -7653 6689 -7601
rect 6701 -7653 6753 -7601
rect 6765 -7653 6817 -7601
rect 6829 -7653 6881 -7601
rect 7281 -7663 7333 -7611
rect 7905 -7649 7957 -7597
rect 7969 -7649 8021 -7597
rect 8033 -7649 8085 -7597
rect 8097 -7649 8149 -7597
rect 8545 -7657 8597 -7605
rect 3778 -8156 3830 -8104
rect 3842 -8156 3894 -8104
rect 3906 -8156 3958 -8104
rect 3970 -8156 4022 -8104
rect 4034 -8156 4086 -8104
rect 4098 -8156 4150 -8104
rect 4162 -8156 4214 -8104
rect 4226 -8156 4278 -8104
rect 4290 -8156 4342 -8104
rect 4354 -8156 4406 -8104
rect 4418 -8156 4470 -8104
rect 4482 -8156 4534 -8104
rect 4546 -8156 4598 -8104
rect 4610 -8156 4662 -8104
rect 4674 -8156 4726 -8104
rect 5020 -8156 5072 -8104
rect 5084 -8156 5136 -8104
rect 5148 -8156 5200 -8104
rect 5212 -8156 5264 -8104
rect 5276 -8156 5328 -8104
rect 5340 -8156 5392 -8104
rect 5404 -8156 5456 -8104
rect 5468 -8156 5520 -8104
rect 5532 -8156 5584 -8104
rect 5596 -8156 5648 -8104
rect 5660 -8156 5712 -8104
rect 5724 -8156 5776 -8104
rect 5788 -8156 5840 -8104
rect 5852 -8156 5904 -8104
rect 5916 -8156 5968 -8104
rect 6259 -8150 6311 -8098
rect 6323 -8150 6375 -8098
rect 6387 -8150 6439 -8098
rect 6451 -8150 6503 -8098
rect 6515 -8150 6567 -8098
rect 6579 -8150 6631 -8098
rect 6643 -8150 6695 -8098
rect 6707 -8150 6759 -8098
rect 6771 -8150 6823 -8098
rect 6835 -8150 6887 -8098
rect 6899 -8150 6951 -8098
rect 6963 -8150 7015 -8098
rect 7027 -8150 7079 -8098
rect 7091 -8150 7143 -8098
rect 7155 -8150 7207 -8098
rect 7521 -8155 7573 -8103
rect 7585 -8155 7637 -8103
rect 7649 -8155 7701 -8103
rect 7713 -8155 7765 -8103
rect 7777 -8155 7829 -8103
rect 7841 -8155 7893 -8103
rect 7905 -8155 7957 -8103
rect 7969 -8155 8021 -8103
rect 8033 -8155 8085 -8103
rect 8097 -8155 8149 -8103
rect 8161 -8155 8213 -8103
rect 8225 -8155 8277 -8103
rect 8289 -8155 8341 -8103
rect 8353 -8155 8405 -8103
rect 8417 -8155 8469 -8103
rect 9604 -8156 9656 -8104
<< metal2 >>
rect 1890 281 10700 300
rect 1890 276 3628 281
rect 1890 224 1914 276
rect 1966 229 3628 276
rect 3680 229 3692 281
rect 3744 229 3756 281
rect 3808 229 3820 281
rect 3872 271 7824 281
rect 3872 229 6240 271
rect 1966 224 6240 229
rect 1890 219 6240 224
rect 6292 229 7824 271
rect 7876 229 7888 281
rect 7940 229 7952 281
rect 8004 229 8016 281
rect 8068 278 10700 281
rect 8068 229 10539 278
rect 6292 226 10539 229
rect 10591 226 10700 278
rect 6292 219 10700 226
rect 1890 200 10700 219
rect 6540 128 10420 140
rect 6540 72 6562 128
rect 6618 72 10352 128
rect 10408 72 10420 128
rect 6540 60 10420 72
rect 7640 -332 7720 -310
rect 7640 -388 7652 -332
rect 7708 -388 7720 -332
rect 7640 -412 7720 -388
rect 7640 -468 7652 -412
rect 7708 -468 7720 -412
rect 7640 -490 7720 -468
rect 2030 -540 2108 -537
rect 2020 -553 12800 -540
rect 2020 -605 2043 -553
rect 2095 -605 2951 -553
rect 3003 -605 3015 -553
rect 3067 -605 3079 -553
rect 3131 -605 3143 -553
rect 3195 -605 3207 -553
rect 3259 -605 3271 -553
rect 3323 -605 3335 -553
rect 3387 -605 3399 -553
rect 3451 -605 3463 -553
rect 3515 -605 3527 -553
rect 3579 -605 3591 -553
rect 3643 -605 3655 -553
rect 3707 -605 3719 -553
rect 3771 -605 3783 -553
rect 3835 -605 3847 -553
rect 3899 -555 12800 -553
rect 3899 -557 5474 -555
rect 3899 -605 4210 -557
rect 2020 -609 4210 -605
rect 4262 -609 4274 -557
rect 4326 -609 4338 -557
rect 4390 -609 4402 -557
rect 4454 -609 4466 -557
rect 4518 -609 4530 -557
rect 4582 -609 4594 -557
rect 4646 -609 4658 -557
rect 4710 -609 4722 -557
rect 4774 -609 4786 -557
rect 4838 -609 4850 -557
rect 4902 -609 4914 -557
rect 4966 -609 4978 -557
rect 5030 -609 5042 -557
rect 5094 -609 5106 -557
rect 5158 -607 5474 -557
rect 5526 -607 5538 -555
rect 5590 -607 5602 -555
rect 5654 -607 5666 -555
rect 5718 -607 5730 -555
rect 5782 -607 5794 -555
rect 5846 -607 5858 -555
rect 5910 -607 5922 -555
rect 5974 -607 5986 -555
rect 6038 -607 6050 -555
rect 6102 -607 6114 -555
rect 6166 -607 6178 -555
rect 6230 -607 6242 -555
rect 6294 -607 6306 -555
rect 6358 -607 6370 -555
rect 6422 -557 12800 -555
rect 6422 -559 7993 -557
rect 6422 -607 6738 -559
rect 5158 -609 6738 -607
rect 2020 -611 6738 -609
rect 6790 -611 6802 -559
rect 6854 -611 6866 -559
rect 6918 -611 6930 -559
rect 6982 -611 6994 -559
rect 7046 -611 7058 -559
rect 7110 -611 7122 -559
rect 7174 -611 7186 -559
rect 7238 -611 7250 -559
rect 7302 -611 7314 -559
rect 7366 -611 7378 -559
rect 7430 -611 7442 -559
rect 7494 -611 7506 -559
rect 7558 -611 7570 -559
rect 7622 -611 7634 -559
rect 7686 -609 7993 -559
rect 8045 -609 8057 -557
rect 8109 -609 8121 -557
rect 8173 -609 8185 -557
rect 8237 -609 8249 -557
rect 8301 -609 8313 -557
rect 8365 -609 8377 -557
rect 8429 -609 8441 -557
rect 8493 -609 8505 -557
rect 8557 -609 8569 -557
rect 8621 -609 8633 -557
rect 8685 -609 8697 -557
rect 8749 -609 8761 -557
rect 8813 -609 8825 -557
rect 8877 -609 8889 -557
rect 8941 -609 9264 -557
rect 9316 -609 9328 -557
rect 9380 -609 9392 -557
rect 9444 -609 9456 -557
rect 9508 -609 9520 -557
rect 9572 -609 9584 -557
rect 9636 -609 9648 -557
rect 9700 -609 9712 -557
rect 9764 -609 9776 -557
rect 9828 -609 9840 -557
rect 9892 -609 9904 -557
rect 9956 -609 9968 -557
rect 10020 -609 10032 -557
rect 10084 -609 10096 -557
rect 10148 -609 10160 -557
rect 10212 -560 12800 -557
rect 10212 -609 10527 -560
rect 7686 -611 10527 -609
rect 2020 -612 10527 -611
rect 10579 -612 10591 -560
rect 10643 -612 10655 -560
rect 10707 -612 10719 -560
rect 10771 -612 10783 -560
rect 10835 -612 10847 -560
rect 10899 -612 10911 -560
rect 10963 -612 10975 -560
rect 11027 -612 11039 -560
rect 11091 -612 11103 -560
rect 11155 -612 11167 -560
rect 11219 -612 11231 -560
rect 11283 -612 11295 -560
rect 11347 -612 11359 -560
rect 11411 -612 11423 -560
rect 11475 -612 11790 -560
rect 11842 -612 11854 -560
rect 11906 -612 11918 -560
rect 11970 -612 11982 -560
rect 12034 -612 12046 -560
rect 12098 -612 12110 -560
rect 12162 -612 12174 -560
rect 12226 -612 12238 -560
rect 12290 -612 12302 -560
rect 12354 -612 12366 -560
rect 12418 -612 12430 -560
rect 12482 -612 12494 -560
rect 12546 -612 12558 -560
rect 12610 -612 12622 -560
rect 12674 -612 12686 -560
rect 12738 -612 12800 -560
rect 2020 -620 12800 -612
rect 2030 -621 2108 -620
rect 6560 -682 6620 -670
rect 3980 -752 4060 -730
rect 3980 -808 3992 -752
rect 4048 -808 4060 -752
rect 3980 -814 3994 -808
rect 4046 -814 4060 -808
rect 3980 -826 4060 -814
rect 3980 -832 3994 -826
rect 4046 -832 4060 -826
rect 3980 -888 3992 -832
rect 4048 -888 4060 -832
rect 3980 -910 4060 -888
rect 5240 -752 5320 -730
rect 5240 -808 5252 -752
rect 5308 -808 5320 -752
rect 5240 -814 5254 -808
rect 5306 -814 5320 -808
rect 5240 -826 5320 -814
rect 5240 -832 5254 -826
rect 5306 -832 5320 -826
rect 5240 -888 5252 -832
rect 5308 -888 5320 -832
rect 5240 -910 5320 -888
rect 6560 -738 6562 -682
rect 6618 -738 6620 -682
rect 10352 -724 10412 -695
rect 6560 -760 6564 -738
rect 6616 -760 6620 -738
rect 6560 -762 6620 -760
rect 6560 -818 6562 -762
rect 6618 -818 6620 -762
rect 6560 -824 6564 -818
rect 6616 -824 6620 -818
rect 6560 -836 6620 -824
rect 6560 -842 6564 -836
rect 6616 -842 6620 -836
rect 6560 -898 6562 -842
rect 6618 -898 6620 -842
rect 6560 -900 6620 -898
rect 6560 -922 6564 -900
rect 6616 -922 6620 -900
rect 7760 -752 7840 -730
rect 7760 -808 7772 -752
rect 7828 -808 7840 -752
rect 7760 -814 7774 -808
rect 7826 -814 7840 -808
rect 7760 -826 7840 -814
rect 7760 -832 7774 -826
rect 7826 -832 7840 -826
rect 7760 -888 7772 -832
rect 7828 -888 7840 -832
rect 7760 -910 7840 -888
rect 9020 -752 9100 -730
rect 9020 -808 9032 -752
rect 9088 -808 9100 -752
rect 9020 -814 9034 -808
rect 9086 -814 9100 -808
rect 9020 -826 9100 -814
rect 9020 -832 9034 -826
rect 9086 -832 9100 -826
rect 9020 -888 9032 -832
rect 9088 -888 9100 -832
rect 9020 -910 9100 -888
rect 10352 -738 10356 -724
rect 10408 -738 10412 -724
rect 10352 -794 10354 -738
rect 10410 -794 10412 -738
rect 10352 -818 10356 -794
rect 10408 -818 10412 -794
rect 10352 -874 10354 -818
rect 10410 -874 10412 -818
rect 10352 -898 10356 -874
rect 10408 -898 10412 -874
rect 6560 -978 6562 -922
rect 6618 -978 6620 -922
rect 6560 -990 6620 -978
rect 10352 -954 10354 -898
rect 10410 -954 10412 -898
rect 11560 -752 11640 -730
rect 11560 -808 11572 -752
rect 11628 -808 11640 -752
rect 11560 -814 11574 -808
rect 11626 -814 11640 -808
rect 11560 -826 11640 -814
rect 11560 -832 11574 -826
rect 11626 -832 11640 -826
rect 11560 -888 11572 -832
rect 11628 -888 11640 -832
rect 11560 -910 11640 -888
rect 12820 -752 12900 -730
rect 12820 -808 12832 -752
rect 12888 -808 12900 -752
rect 12820 -814 12834 -808
rect 12886 -814 12900 -808
rect 12820 -826 12900 -814
rect 12820 -832 12834 -826
rect 12886 -832 12900 -826
rect 12820 -888 12832 -832
rect 12888 -888 12900 -832
rect 12820 -910 12900 -888
rect 10352 -968 10356 -954
rect 10408 -968 10412 -954
rect 10352 -996 10412 -968
rect 9250 -1020 10233 -1018
rect 2159 -1040 2218 -1038
rect 2700 -1040 5189 -1030
rect 2150 -1048 5189 -1040
rect 5271 -1042 5332 -1036
rect 5472 -1038 6438 -1027
rect 9240 -1034 10240 -1020
rect 5472 -1040 5481 -1038
rect 2150 -1055 2993 -1048
rect 2150 -1107 2162 -1055
rect 2214 -1100 2993 -1055
rect 3045 -1100 3057 -1048
rect 3109 -1100 3121 -1048
rect 3173 -1100 3185 -1048
rect 3237 -1100 3249 -1048
rect 3301 -1100 3313 -1048
rect 3365 -1100 3377 -1048
rect 3429 -1100 3441 -1048
rect 3493 -1100 3505 -1048
rect 3557 -1100 3569 -1048
rect 3621 -1100 3633 -1048
rect 3685 -1100 3697 -1048
rect 3749 -1100 3761 -1048
rect 3813 -1100 3825 -1048
rect 3877 -1050 5189 -1048
rect 3877 -1100 4239 -1050
rect 2214 -1102 4239 -1100
rect 4291 -1102 4303 -1050
rect 4355 -1102 4367 -1050
rect 4419 -1102 4431 -1050
rect 4483 -1102 4495 -1050
rect 4547 -1102 4559 -1050
rect 4611 -1102 4623 -1050
rect 4675 -1102 4687 -1050
rect 4739 -1102 4751 -1050
rect 4803 -1102 4815 -1050
rect 4867 -1102 4879 -1050
rect 4931 -1102 4943 -1050
rect 4995 -1102 5007 -1050
rect 5059 -1102 5071 -1050
rect 5123 -1102 5189 -1050
rect 2214 -1107 5189 -1102
rect 2150 -1120 5189 -1107
rect 5260 -1054 5337 -1042
rect 5260 -1106 5275 -1054
rect 5327 -1060 5337 -1054
rect 5440 -1060 5481 -1040
rect 5327 -1090 5481 -1060
rect 5533 -1090 5545 -1038
rect 5597 -1090 5609 -1038
rect 5661 -1090 5673 -1038
rect 5725 -1090 5737 -1038
rect 5789 -1090 5801 -1038
rect 5853 -1090 5865 -1038
rect 5917 -1090 5929 -1038
rect 5981 -1090 5993 -1038
rect 6045 -1090 6057 -1038
rect 6109 -1090 6121 -1038
rect 6173 -1090 6185 -1038
rect 6237 -1090 6249 -1038
rect 6301 -1090 6313 -1038
rect 6365 -1090 6377 -1038
rect 6429 -1040 6438 -1038
rect 6429 -1090 6460 -1040
rect 5327 -1106 6460 -1090
rect 5260 -1120 6460 -1106
rect 6700 -1046 8960 -1040
rect 9050 -1041 9109 -1038
rect 6700 -1098 6746 -1046
rect 6798 -1098 6810 -1046
rect 6862 -1098 6874 -1046
rect 6926 -1098 6938 -1046
rect 6990 -1098 7002 -1046
rect 7054 -1098 7066 -1046
rect 7118 -1098 7130 -1046
rect 7182 -1098 7194 -1046
rect 7246 -1098 7258 -1046
rect 7310 -1098 7322 -1046
rect 7374 -1098 7386 -1046
rect 7438 -1098 7450 -1046
rect 7502 -1098 7514 -1046
rect 7566 -1098 7578 -1046
rect 7630 -1059 8004 -1046
rect 7630 -1098 7853 -1059
rect 6700 -1115 7853 -1098
rect 7909 -1098 8004 -1059
rect 8056 -1098 8068 -1046
rect 8120 -1098 8132 -1046
rect 8184 -1098 8196 -1046
rect 8248 -1098 8260 -1046
rect 8312 -1098 8324 -1046
rect 8376 -1098 8388 -1046
rect 8440 -1098 8452 -1046
rect 8504 -1098 8516 -1046
rect 8568 -1098 8580 -1046
rect 8632 -1098 8644 -1046
rect 8696 -1098 8708 -1046
rect 8760 -1098 8772 -1046
rect 8824 -1098 8836 -1046
rect 8888 -1098 8960 -1046
rect 9040 -1054 9119 -1041
rect 9040 -1083 9053 -1054
rect 7909 -1115 8960 -1098
rect 6700 -1120 8960 -1115
rect 9041 -1106 9053 -1083
rect 9105 -1061 9119 -1054
rect 9240 -1061 9267 -1034
rect 9105 -1086 9267 -1061
rect 9319 -1086 9331 -1034
rect 9383 -1086 9395 -1034
rect 9447 -1086 9459 -1034
rect 9511 -1086 9523 -1034
rect 9575 -1086 9587 -1034
rect 9639 -1086 9651 -1034
rect 9703 -1086 9715 -1034
rect 9767 -1086 9779 -1034
rect 9831 -1086 9843 -1034
rect 9895 -1086 9907 -1034
rect 9959 -1086 9971 -1034
rect 10023 -1086 10035 -1034
rect 10087 -1086 10099 -1034
rect 10151 -1086 10163 -1034
rect 10215 -1086 10240 -1034
rect 9105 -1100 10240 -1086
rect 10500 -1049 13960 -1030
rect 9105 -1106 10239 -1100
rect 2159 -1123 2218 -1120
rect 5271 -1124 5332 -1120
rect 7832 -1128 7930 -1120
rect 9041 -1125 10239 -1106
rect 10500 -1101 10548 -1049
rect 10600 -1101 10612 -1049
rect 10664 -1101 10676 -1049
rect 10728 -1101 10740 -1049
rect 10792 -1101 10804 -1049
rect 10856 -1101 10868 -1049
rect 10920 -1101 10932 -1049
rect 10984 -1101 10996 -1049
rect 11048 -1101 11060 -1049
rect 11112 -1101 11124 -1049
rect 11176 -1101 11188 -1049
rect 11240 -1101 11252 -1049
rect 11304 -1101 11316 -1049
rect 11368 -1101 11380 -1049
rect 11432 -1052 13960 -1049
rect 11432 -1056 13892 -1052
rect 11432 -1101 11814 -1056
rect 10500 -1108 11814 -1101
rect 11866 -1108 11878 -1056
rect 11930 -1108 11942 -1056
rect 11994 -1108 12006 -1056
rect 12058 -1108 12070 -1056
rect 12122 -1108 12134 -1056
rect 12186 -1108 12198 -1056
rect 12250 -1108 12262 -1056
rect 12314 -1108 12326 -1056
rect 12378 -1108 12390 -1056
rect 12442 -1108 12454 -1056
rect 12506 -1108 12518 -1056
rect 12570 -1108 12582 -1056
rect 12634 -1108 12646 -1056
rect 12698 -1104 13892 -1056
rect 13944 -1104 13960 -1052
rect 12698 -1108 13960 -1104
rect 10500 -1120 13960 -1108
rect 2031 -1220 2109 -1215
rect 2020 -1231 12800 -1220
rect 2020 -1283 2044 -1231
rect 2096 -1236 8020 -1231
rect 2096 -1283 2951 -1236
rect 2020 -1288 2951 -1283
rect 3003 -1288 3015 -1236
rect 3067 -1288 3079 -1236
rect 3131 -1288 3143 -1236
rect 3195 -1288 3207 -1236
rect 3259 -1288 3271 -1236
rect 3323 -1288 3335 -1236
rect 3387 -1288 3399 -1236
rect 3451 -1288 3463 -1236
rect 3515 -1288 3527 -1236
rect 3579 -1288 3591 -1236
rect 3643 -1288 3655 -1236
rect 3707 -1288 3719 -1236
rect 3771 -1288 3783 -1236
rect 3835 -1288 3847 -1236
rect 3899 -1237 8020 -1236
rect 3899 -1242 5498 -1237
rect 3899 -1288 4220 -1242
rect 2020 -1294 4220 -1288
rect 4272 -1294 4284 -1242
rect 4336 -1294 4348 -1242
rect 4400 -1294 4412 -1242
rect 4464 -1294 4476 -1242
rect 4528 -1294 4540 -1242
rect 4592 -1294 4604 -1242
rect 4656 -1294 4668 -1242
rect 4720 -1294 4732 -1242
rect 4784 -1294 4796 -1242
rect 4848 -1294 4860 -1242
rect 4912 -1294 4924 -1242
rect 4976 -1294 4988 -1242
rect 5040 -1294 5052 -1242
rect 5104 -1294 5116 -1242
rect 5168 -1289 5498 -1242
rect 5550 -1289 5562 -1237
rect 5614 -1289 5626 -1237
rect 5678 -1289 5690 -1237
rect 5742 -1289 5754 -1237
rect 5806 -1289 5818 -1237
rect 5870 -1289 5882 -1237
rect 5934 -1289 5946 -1237
rect 5998 -1289 6010 -1237
rect 6062 -1289 6074 -1237
rect 6126 -1289 6138 -1237
rect 6190 -1289 6202 -1237
rect 6254 -1289 6266 -1237
rect 6318 -1289 6330 -1237
rect 6382 -1289 6737 -1237
rect 6789 -1289 6801 -1237
rect 6853 -1289 6865 -1237
rect 6917 -1289 6929 -1237
rect 6981 -1289 6993 -1237
rect 7045 -1289 7057 -1237
rect 7109 -1289 7121 -1237
rect 7173 -1289 7185 -1237
rect 7237 -1289 7249 -1237
rect 7301 -1289 7313 -1237
rect 7365 -1289 7377 -1237
rect 7429 -1289 7441 -1237
rect 7493 -1289 7505 -1237
rect 7557 -1289 7569 -1237
rect 7621 -1289 7633 -1237
rect 7685 -1283 8020 -1237
rect 8072 -1283 8084 -1231
rect 8136 -1283 8148 -1231
rect 8200 -1283 8212 -1231
rect 8264 -1283 8276 -1231
rect 8328 -1283 8340 -1231
rect 8392 -1283 8404 -1231
rect 8456 -1283 8468 -1231
rect 8520 -1283 8532 -1231
rect 8584 -1283 8596 -1231
rect 8648 -1283 8660 -1231
rect 8712 -1283 8724 -1231
rect 8776 -1283 8788 -1231
rect 8840 -1283 8852 -1231
rect 8904 -1237 12800 -1231
rect 8904 -1243 11783 -1237
rect 8904 -1283 9283 -1243
rect 7685 -1289 9283 -1283
rect 5168 -1294 9283 -1289
rect 2020 -1295 9283 -1294
rect 9335 -1295 9347 -1243
rect 9399 -1295 9411 -1243
rect 9463 -1295 9475 -1243
rect 9527 -1295 9539 -1243
rect 9591 -1295 9603 -1243
rect 9655 -1295 9667 -1243
rect 9719 -1295 9731 -1243
rect 9783 -1295 9795 -1243
rect 9847 -1295 9859 -1243
rect 9911 -1295 9923 -1243
rect 9975 -1295 9987 -1243
rect 10039 -1295 10051 -1243
rect 10103 -1295 10115 -1243
rect 10167 -1295 10525 -1243
rect 10577 -1295 10589 -1243
rect 10641 -1295 10653 -1243
rect 10705 -1295 10717 -1243
rect 10769 -1295 10781 -1243
rect 10833 -1295 10845 -1243
rect 10897 -1295 10909 -1243
rect 10961 -1295 10973 -1243
rect 11025 -1295 11037 -1243
rect 11089 -1295 11101 -1243
rect 11153 -1295 11165 -1243
rect 11217 -1295 11229 -1243
rect 11281 -1295 11293 -1243
rect 11345 -1295 11357 -1243
rect 11409 -1295 11421 -1243
rect 11473 -1289 11783 -1243
rect 11835 -1289 11847 -1237
rect 11899 -1289 11911 -1237
rect 11963 -1289 11975 -1237
rect 12027 -1289 12039 -1237
rect 12091 -1289 12103 -1237
rect 12155 -1289 12167 -1237
rect 12219 -1289 12231 -1237
rect 12283 -1289 12295 -1237
rect 12347 -1289 12359 -1237
rect 12411 -1289 12423 -1237
rect 12475 -1289 12487 -1237
rect 12539 -1289 12551 -1237
rect 12603 -1289 12615 -1237
rect 12667 -1289 12679 -1237
rect 12731 -1289 12800 -1237
rect 11473 -1295 12800 -1289
rect 2020 -1300 12800 -1295
rect 3980 -1452 4060 -1430
rect 3980 -1508 3992 -1452
rect 4048 -1508 4060 -1452
rect 3980 -1514 3994 -1508
rect 4046 -1514 4060 -1508
rect 3980 -1526 4060 -1514
rect 3980 -1532 3994 -1526
rect 4046 -1532 4060 -1526
rect 3980 -1588 3992 -1532
rect 4048 -1588 4060 -1532
rect 3980 -1610 4060 -1588
rect 5260 -1452 5340 -1430
rect 5260 -1508 5272 -1452
rect 5328 -1508 5340 -1452
rect 5260 -1514 5274 -1508
rect 5326 -1514 5340 -1508
rect 5260 -1526 5340 -1514
rect 5260 -1532 5274 -1526
rect 5326 -1532 5340 -1526
rect 5260 -1588 5272 -1532
rect 5328 -1588 5340 -1532
rect 5260 -1610 5340 -1588
rect 9040 -1452 9120 -1430
rect 9040 -1508 9052 -1452
rect 9108 -1508 9120 -1452
rect 9040 -1514 9054 -1508
rect 9106 -1514 9120 -1508
rect 9040 -1526 9120 -1514
rect 9040 -1532 9054 -1526
rect 9106 -1532 9120 -1526
rect 9040 -1588 9052 -1532
rect 9108 -1588 9120 -1532
rect 9040 -1610 9120 -1588
rect 11560 -1452 11640 -1430
rect 11560 -1508 11572 -1452
rect 11628 -1508 11640 -1452
rect 11560 -1514 11574 -1508
rect 11626 -1514 11640 -1508
rect 11560 -1526 11640 -1514
rect 11560 -1532 11574 -1526
rect 11626 -1532 11640 -1526
rect 11560 -1588 11572 -1532
rect 11628 -1588 11640 -1532
rect 11560 -1610 11640 -1588
rect 12820 -1452 12900 -1430
rect 12820 -1508 12832 -1452
rect 12888 -1508 12900 -1452
rect 12820 -1514 12834 -1508
rect 12886 -1514 12900 -1508
rect 12820 -1526 12900 -1514
rect 12820 -1532 12834 -1526
rect 12886 -1532 12900 -1526
rect 12820 -1588 12832 -1532
rect 12888 -1588 12900 -1532
rect 12820 -1610 12900 -1588
rect 1780 -1710 1862 -1700
rect 1780 -1727 5189 -1710
rect 6650 -1720 6708 -1719
rect 1780 -1779 1793 -1727
rect 1845 -1732 4243 -1727
rect 1845 -1779 2974 -1732
rect 1780 -1784 2974 -1779
rect 3026 -1784 3038 -1732
rect 3090 -1784 3102 -1732
rect 3154 -1784 3166 -1732
rect 3218 -1784 3230 -1732
rect 3282 -1784 3294 -1732
rect 3346 -1784 3358 -1732
rect 3410 -1784 3422 -1732
rect 3474 -1784 3486 -1732
rect 3538 -1784 3550 -1732
rect 3602 -1784 3614 -1732
rect 3666 -1784 3678 -1732
rect 3730 -1784 3742 -1732
rect 3794 -1784 3806 -1732
rect 3858 -1779 4243 -1732
rect 4295 -1779 4307 -1727
rect 4359 -1779 4371 -1727
rect 4423 -1779 4435 -1727
rect 4487 -1779 4499 -1727
rect 4551 -1779 4563 -1727
rect 4615 -1779 4627 -1727
rect 4679 -1779 4691 -1727
rect 4743 -1779 4755 -1727
rect 4807 -1779 4819 -1727
rect 4871 -1779 4883 -1727
rect 4935 -1779 4947 -1727
rect 4999 -1779 5011 -1727
rect 5063 -1779 5075 -1727
rect 5127 -1779 5189 -1727
rect 3858 -1784 5189 -1779
rect 1780 -1800 5189 -1784
rect 6623 -1734 8980 -1720
rect 6623 -1737 8021 -1734
rect 6623 -1753 6762 -1737
rect 6623 -1809 6649 -1753
rect 6705 -1789 6762 -1753
rect 6814 -1789 6826 -1737
rect 6878 -1789 6890 -1737
rect 6942 -1789 6954 -1737
rect 7006 -1789 7018 -1737
rect 7070 -1789 7082 -1737
rect 7134 -1789 7146 -1737
rect 7198 -1789 7210 -1737
rect 7262 -1789 7274 -1737
rect 7326 -1789 7338 -1737
rect 7390 -1789 7402 -1737
rect 7454 -1789 7466 -1737
rect 7518 -1789 7530 -1737
rect 7582 -1789 7594 -1737
rect 7646 -1786 8021 -1737
rect 8073 -1786 8085 -1734
rect 8137 -1786 8149 -1734
rect 8201 -1786 8213 -1734
rect 8265 -1786 8277 -1734
rect 8329 -1786 8341 -1734
rect 8393 -1786 8405 -1734
rect 8457 -1786 8469 -1734
rect 8521 -1786 8533 -1734
rect 8585 -1786 8597 -1734
rect 8649 -1786 8661 -1734
rect 8713 -1786 8725 -1734
rect 8777 -1786 8789 -1734
rect 8841 -1786 8853 -1734
rect 8905 -1786 8980 -1734
rect 7646 -1789 8980 -1786
rect 6705 -1800 8980 -1789
rect 10500 -1726 13850 -1710
rect 10500 -1727 13782 -1726
rect 10500 -1779 10566 -1727
rect 10618 -1779 10630 -1727
rect 10682 -1779 10694 -1727
rect 10746 -1779 10758 -1727
rect 10810 -1779 10822 -1727
rect 10874 -1779 10886 -1727
rect 10938 -1779 10950 -1727
rect 11002 -1779 11014 -1727
rect 11066 -1779 11078 -1727
rect 11130 -1779 11142 -1727
rect 11194 -1779 11206 -1727
rect 11258 -1779 11270 -1727
rect 11322 -1779 11334 -1727
rect 11386 -1779 11398 -1727
rect 11450 -1732 13782 -1727
rect 11450 -1779 11812 -1732
rect 10500 -1784 11812 -1779
rect 11864 -1784 11876 -1732
rect 11928 -1784 11940 -1732
rect 11992 -1784 12004 -1732
rect 12056 -1784 12068 -1732
rect 12120 -1784 12132 -1732
rect 12184 -1784 12196 -1732
rect 12248 -1784 12260 -1732
rect 12312 -1784 12324 -1732
rect 12376 -1784 12388 -1732
rect 12440 -1784 12452 -1732
rect 12504 -1784 12516 -1732
rect 12568 -1784 12580 -1732
rect 12632 -1784 12644 -1732
rect 12696 -1778 13782 -1732
rect 13834 -1778 13850 -1726
rect 12696 -1784 13850 -1778
rect 10500 -1800 13850 -1784
rect 6705 -1809 6716 -1800
rect 6623 -1834 6716 -1809
rect 6647 -1839 6708 -1834
rect 2031 -1900 2109 -1899
rect 2020 -1911 12820 -1900
rect 2020 -1915 2950 -1911
rect 2020 -1967 2044 -1915
rect 2096 -1963 2950 -1915
rect 3002 -1963 3014 -1911
rect 3066 -1963 3078 -1911
rect 3130 -1963 3142 -1911
rect 3194 -1963 3206 -1911
rect 3258 -1963 3270 -1911
rect 3322 -1963 3334 -1911
rect 3386 -1963 3398 -1911
rect 3450 -1963 3462 -1911
rect 3514 -1963 3526 -1911
rect 3578 -1963 3590 -1911
rect 3642 -1963 3654 -1911
rect 3706 -1963 3718 -1911
rect 3770 -1963 3782 -1911
rect 3834 -1963 3846 -1911
rect 3898 -1913 12820 -1911
rect 3898 -1921 5480 -1913
rect 3898 -1963 4216 -1921
rect 2096 -1967 4216 -1963
rect 2020 -1973 4216 -1967
rect 4268 -1973 4280 -1921
rect 4332 -1973 4344 -1921
rect 4396 -1973 4408 -1921
rect 4460 -1973 4472 -1921
rect 4524 -1973 4536 -1921
rect 4588 -1973 4600 -1921
rect 4652 -1973 4664 -1921
rect 4716 -1973 4728 -1921
rect 4780 -1973 4792 -1921
rect 4844 -1973 4856 -1921
rect 4908 -1973 4920 -1921
rect 4972 -1973 4984 -1921
rect 5036 -1973 5048 -1921
rect 5100 -1973 5112 -1921
rect 5164 -1965 5480 -1921
rect 5532 -1965 5544 -1913
rect 5596 -1965 5608 -1913
rect 5660 -1965 5672 -1913
rect 5724 -1965 5736 -1913
rect 5788 -1965 5800 -1913
rect 5852 -1965 5864 -1913
rect 5916 -1965 5928 -1913
rect 5980 -1965 5992 -1913
rect 6044 -1965 6056 -1913
rect 6108 -1965 6120 -1913
rect 6172 -1965 6184 -1913
rect 6236 -1965 6248 -1913
rect 6300 -1965 6312 -1913
rect 6364 -1965 6376 -1913
rect 6428 -1920 12820 -1913
rect 6428 -1922 9259 -1920
rect 6428 -1965 6739 -1922
rect 5164 -1973 6739 -1965
rect 2020 -1974 6739 -1973
rect 6791 -1974 6803 -1922
rect 6855 -1974 6867 -1922
rect 6919 -1974 6931 -1922
rect 6983 -1974 6995 -1922
rect 7047 -1974 7059 -1922
rect 7111 -1974 7123 -1922
rect 7175 -1974 7187 -1922
rect 7239 -1974 7251 -1922
rect 7303 -1974 7315 -1922
rect 7367 -1974 7379 -1922
rect 7431 -1974 7443 -1922
rect 7495 -1974 7507 -1922
rect 7559 -1974 7571 -1922
rect 7623 -1974 7635 -1922
rect 7687 -1923 9259 -1922
rect 7687 -1974 8000 -1923
rect 2020 -1975 8000 -1974
rect 8052 -1975 8064 -1923
rect 8116 -1975 8128 -1923
rect 8180 -1975 8192 -1923
rect 8244 -1975 8256 -1923
rect 8308 -1975 8320 -1923
rect 8372 -1975 8384 -1923
rect 8436 -1975 8448 -1923
rect 8500 -1975 8512 -1923
rect 8564 -1975 8576 -1923
rect 8628 -1975 8640 -1923
rect 8692 -1975 8704 -1923
rect 8756 -1975 8768 -1923
rect 8820 -1975 8832 -1923
rect 8884 -1975 8896 -1923
rect 8948 -1972 9259 -1923
rect 9311 -1972 9323 -1920
rect 9375 -1972 9387 -1920
rect 9439 -1972 9451 -1920
rect 9503 -1972 9515 -1920
rect 9567 -1972 9579 -1920
rect 9631 -1972 9643 -1920
rect 9695 -1972 9707 -1920
rect 9759 -1972 9771 -1920
rect 9823 -1972 9835 -1920
rect 9887 -1972 9899 -1920
rect 9951 -1972 9963 -1920
rect 10015 -1972 10027 -1920
rect 10079 -1972 10091 -1920
rect 10143 -1972 10155 -1920
rect 10207 -1921 12820 -1920
rect 10207 -1924 11780 -1921
rect 10207 -1972 10521 -1924
rect 8948 -1975 10521 -1972
rect 2020 -1976 10521 -1975
rect 10573 -1976 10585 -1924
rect 10637 -1976 10649 -1924
rect 10701 -1976 10713 -1924
rect 10765 -1976 10777 -1924
rect 10829 -1976 10841 -1924
rect 10893 -1976 10905 -1924
rect 10957 -1976 10969 -1924
rect 11021 -1976 11033 -1924
rect 11085 -1976 11097 -1924
rect 11149 -1976 11161 -1924
rect 11213 -1976 11225 -1924
rect 11277 -1976 11289 -1924
rect 11341 -1976 11353 -1924
rect 11405 -1976 11417 -1924
rect 11469 -1973 11780 -1924
rect 11832 -1973 11844 -1921
rect 11896 -1973 11908 -1921
rect 11960 -1973 11972 -1921
rect 12024 -1973 12036 -1921
rect 12088 -1973 12100 -1921
rect 12152 -1973 12164 -1921
rect 12216 -1973 12228 -1921
rect 12280 -1973 12292 -1921
rect 12344 -1973 12356 -1921
rect 12408 -1973 12420 -1921
rect 12472 -1973 12484 -1921
rect 12536 -1973 12548 -1921
rect 12600 -1973 12612 -1921
rect 12664 -1973 12676 -1921
rect 12728 -1973 12820 -1921
rect 11469 -1976 12820 -1973
rect 2020 -1980 12820 -1976
rect 2031 -1983 2109 -1980
rect 3980 -2152 4060 -2130
rect 3980 -2208 3992 -2152
rect 4048 -2208 4060 -2152
rect 3980 -2214 3994 -2208
rect 4046 -2214 4060 -2208
rect 3980 -2226 4060 -2214
rect 3980 -2232 3994 -2226
rect 4046 -2232 4060 -2226
rect 3980 -2288 3992 -2232
rect 4048 -2288 4060 -2232
rect 3980 -2310 4060 -2288
rect 5240 -2152 5320 -2130
rect 5240 -2208 5252 -2152
rect 5308 -2208 5320 -2152
rect 5240 -2214 5254 -2208
rect 5306 -2214 5320 -2208
rect 5240 -2226 5320 -2214
rect 5240 -2232 5254 -2226
rect 5306 -2232 5320 -2226
rect 5240 -2288 5252 -2232
rect 5308 -2288 5320 -2232
rect 5240 -2310 5320 -2288
rect 9040 -2152 9120 -2130
rect 9040 -2208 9052 -2152
rect 9108 -2208 9120 -2152
rect 9040 -2214 9054 -2208
rect 9106 -2214 9120 -2208
rect 9040 -2226 9120 -2214
rect 9040 -2232 9054 -2226
rect 9106 -2232 9120 -2226
rect 9040 -2288 9052 -2232
rect 9108 -2288 9120 -2232
rect 9040 -2310 9120 -2288
rect 11560 -2152 11640 -2130
rect 11560 -2208 11572 -2152
rect 11628 -2208 11640 -2152
rect 11560 -2214 11574 -2208
rect 11626 -2214 11640 -2208
rect 11560 -2226 11640 -2214
rect 11560 -2232 11574 -2226
rect 11626 -2232 11640 -2226
rect 11560 -2288 11572 -2232
rect 11628 -2288 11640 -2232
rect 11560 -2310 11640 -2288
rect 12820 -2152 12900 -2130
rect 12820 -2208 12832 -2152
rect 12888 -2208 12900 -2152
rect 12820 -2214 12834 -2208
rect 12886 -2214 12900 -2208
rect 12820 -2226 12900 -2214
rect 12820 -2232 12834 -2226
rect 12886 -2232 12900 -2226
rect 12820 -2288 12832 -2232
rect 12888 -2288 12900 -2232
rect 12820 -2310 12900 -2288
rect 6656 -2400 6757 -2398
rect 1670 -2410 1890 -2400
rect 6656 -2403 9000 -2400
rect 6649 -2404 9000 -2403
rect 6643 -2406 9000 -2404
rect 1670 -2420 5189 -2410
rect 1670 -2425 4250 -2420
rect 1670 -2477 1682 -2425
rect 1734 -2477 2974 -2425
rect 3026 -2477 3038 -2425
rect 3090 -2477 3102 -2425
rect 3154 -2477 3166 -2425
rect 3218 -2477 3230 -2425
rect 3282 -2477 3294 -2425
rect 3346 -2477 3358 -2425
rect 3410 -2477 3422 -2425
rect 3474 -2477 3486 -2425
rect 3538 -2477 3550 -2425
rect 3602 -2477 3614 -2425
rect 3666 -2477 3678 -2425
rect 3730 -2477 3742 -2425
rect 3794 -2477 3806 -2425
rect 3858 -2472 4250 -2425
rect 4302 -2472 4314 -2420
rect 4366 -2472 4378 -2420
rect 4430 -2472 4442 -2420
rect 4494 -2472 4506 -2420
rect 4558 -2472 4570 -2420
rect 4622 -2472 4634 -2420
rect 4686 -2472 4698 -2420
rect 4750 -2472 4762 -2420
rect 4814 -2472 4826 -2420
rect 4878 -2472 4890 -2420
rect 4942 -2472 4954 -2420
rect 5006 -2472 5018 -2420
rect 5070 -2472 5082 -2420
rect 5134 -2472 5189 -2420
rect 3858 -2477 5189 -2472
rect 1670 -2500 5189 -2477
rect 6643 -2415 8009 -2406
rect 6643 -2434 6759 -2415
rect 6643 -2490 6651 -2434
rect 6707 -2467 6759 -2434
rect 6811 -2467 6823 -2415
rect 6875 -2467 6887 -2415
rect 6939 -2467 6951 -2415
rect 7003 -2467 7015 -2415
rect 7067 -2467 7079 -2415
rect 7131 -2467 7143 -2415
rect 7195 -2467 7207 -2415
rect 7259 -2467 7271 -2415
rect 7323 -2467 7335 -2415
rect 7387 -2467 7399 -2415
rect 7451 -2467 7463 -2415
rect 7515 -2467 7527 -2415
rect 7579 -2467 7591 -2415
rect 7643 -2458 8009 -2415
rect 8061 -2458 8073 -2406
rect 8125 -2458 8137 -2406
rect 8189 -2458 8201 -2406
rect 8253 -2458 8265 -2406
rect 8317 -2458 8329 -2406
rect 8381 -2458 8393 -2406
rect 8445 -2458 8457 -2406
rect 8509 -2458 8521 -2406
rect 8573 -2458 8585 -2406
rect 8637 -2458 8649 -2406
rect 8701 -2458 8713 -2406
rect 8765 -2458 8777 -2406
rect 8829 -2458 8841 -2406
rect 8893 -2458 9000 -2406
rect 7643 -2467 9000 -2458
rect 6707 -2480 9000 -2467
rect 10500 -2424 13740 -2410
rect 10500 -2476 10564 -2424
rect 10616 -2476 10628 -2424
rect 10680 -2476 10692 -2424
rect 10744 -2476 10756 -2424
rect 10808 -2476 10820 -2424
rect 10872 -2476 10884 -2424
rect 10936 -2476 10948 -2424
rect 11000 -2476 11012 -2424
rect 11064 -2476 11076 -2424
rect 11128 -2476 11140 -2424
rect 11192 -2476 11204 -2424
rect 11256 -2476 11268 -2424
rect 11320 -2476 11332 -2424
rect 11384 -2476 11396 -2424
rect 11448 -2429 13740 -2424
rect 11448 -2476 11812 -2429
rect 6707 -2487 6757 -2480
rect 10500 -2481 11812 -2476
rect 11864 -2481 11876 -2429
rect 11928 -2481 11940 -2429
rect 11992 -2481 12004 -2429
rect 12056 -2481 12068 -2429
rect 12120 -2481 12132 -2429
rect 12184 -2481 12196 -2429
rect 12248 -2481 12260 -2429
rect 12312 -2481 12324 -2429
rect 12376 -2481 12388 -2429
rect 12440 -2481 12452 -2429
rect 12504 -2481 12516 -2429
rect 12568 -2481 12580 -2429
rect 12632 -2481 12644 -2429
rect 12696 -2434 13740 -2429
rect 12696 -2481 13672 -2434
rect 10500 -2486 13672 -2481
rect 13724 -2486 13740 -2434
rect 6707 -2490 6736 -2487
rect 6643 -2518 6736 -2490
rect 10500 -2500 13740 -2486
rect 6649 -2520 6710 -2518
rect 2020 -2612 12820 -2600
rect 2020 -2616 2947 -2612
rect 2020 -2668 2045 -2616
rect 2097 -2664 2947 -2616
rect 2999 -2664 3011 -2612
rect 3063 -2664 3075 -2612
rect 3127 -2664 3139 -2612
rect 3191 -2664 3203 -2612
rect 3255 -2664 3267 -2612
rect 3319 -2664 3331 -2612
rect 3383 -2664 3395 -2612
rect 3447 -2664 3459 -2612
rect 3511 -2664 3523 -2612
rect 3575 -2664 3587 -2612
rect 3639 -2664 3651 -2612
rect 3703 -2664 3715 -2612
rect 3767 -2664 3779 -2612
rect 3831 -2664 3843 -2612
rect 3895 -2616 12820 -2612
rect 3895 -2617 10525 -2616
rect 3895 -2620 9264 -2617
rect 3895 -2664 4213 -2620
rect 2097 -2668 4213 -2664
rect 2020 -2672 4213 -2668
rect 4265 -2672 4277 -2620
rect 4329 -2672 4341 -2620
rect 4393 -2672 4405 -2620
rect 4457 -2672 4469 -2620
rect 4521 -2672 4533 -2620
rect 4585 -2672 4597 -2620
rect 4649 -2672 4661 -2620
rect 4713 -2672 4725 -2620
rect 4777 -2672 4789 -2620
rect 4841 -2672 4853 -2620
rect 4905 -2672 4917 -2620
rect 4969 -2672 4981 -2620
rect 5033 -2672 5045 -2620
rect 5097 -2672 5109 -2620
rect 5161 -2672 5479 -2620
rect 5531 -2672 5543 -2620
rect 5595 -2672 5607 -2620
rect 5659 -2672 5671 -2620
rect 5723 -2672 5735 -2620
rect 5787 -2672 5799 -2620
rect 5851 -2672 5863 -2620
rect 5915 -2672 5927 -2620
rect 5979 -2672 5991 -2620
rect 6043 -2672 6055 -2620
rect 6107 -2672 6119 -2620
rect 6171 -2672 6183 -2620
rect 6235 -2672 6247 -2620
rect 6299 -2672 6311 -2620
rect 6363 -2672 6375 -2620
rect 6427 -2672 6736 -2620
rect 6788 -2672 6800 -2620
rect 6852 -2672 6864 -2620
rect 6916 -2672 6928 -2620
rect 6980 -2672 6992 -2620
rect 7044 -2672 7056 -2620
rect 7108 -2672 7120 -2620
rect 7172 -2672 7184 -2620
rect 7236 -2672 7248 -2620
rect 7300 -2672 7312 -2620
rect 7364 -2672 7376 -2620
rect 7428 -2672 7440 -2620
rect 7492 -2672 7504 -2620
rect 7556 -2672 7568 -2620
rect 7620 -2672 7632 -2620
rect 7684 -2672 8004 -2620
rect 8056 -2672 8068 -2620
rect 8120 -2672 8132 -2620
rect 8184 -2672 8196 -2620
rect 8248 -2672 8260 -2620
rect 8312 -2672 8324 -2620
rect 8376 -2672 8388 -2620
rect 8440 -2672 8452 -2620
rect 8504 -2672 8516 -2620
rect 8568 -2672 8580 -2620
rect 8632 -2672 8644 -2620
rect 8696 -2672 8708 -2620
rect 8760 -2672 8772 -2620
rect 8824 -2672 8836 -2620
rect 8888 -2672 8900 -2620
rect 8952 -2669 9264 -2620
rect 9316 -2669 9328 -2617
rect 9380 -2669 9392 -2617
rect 9444 -2669 9456 -2617
rect 9508 -2669 9520 -2617
rect 9572 -2669 9584 -2617
rect 9636 -2669 9648 -2617
rect 9700 -2669 9712 -2617
rect 9764 -2669 9776 -2617
rect 9828 -2669 9840 -2617
rect 9892 -2669 9904 -2617
rect 9956 -2669 9968 -2617
rect 10020 -2669 10032 -2617
rect 10084 -2669 10096 -2617
rect 10148 -2669 10160 -2617
rect 10212 -2668 10525 -2617
rect 10577 -2668 10589 -2616
rect 10641 -2668 10653 -2616
rect 10705 -2668 10717 -2616
rect 10769 -2668 10781 -2616
rect 10833 -2668 10845 -2616
rect 10897 -2668 10909 -2616
rect 10961 -2668 10973 -2616
rect 11025 -2668 11037 -2616
rect 11089 -2668 11101 -2616
rect 11153 -2668 11165 -2616
rect 11217 -2668 11229 -2616
rect 11281 -2668 11293 -2616
rect 11345 -2668 11357 -2616
rect 11409 -2668 11421 -2616
rect 11473 -2621 12820 -2616
rect 11473 -2668 11789 -2621
rect 10212 -2669 11789 -2668
rect 8952 -2672 11789 -2669
rect 2020 -2673 11789 -2672
rect 11841 -2673 11853 -2621
rect 11905 -2673 11917 -2621
rect 11969 -2673 11981 -2621
rect 12033 -2673 12045 -2621
rect 12097 -2673 12109 -2621
rect 12161 -2673 12173 -2621
rect 12225 -2673 12237 -2621
rect 12289 -2673 12301 -2621
rect 12353 -2673 12365 -2621
rect 12417 -2673 12429 -2621
rect 12481 -2673 12493 -2621
rect 12545 -2673 12557 -2621
rect 12609 -2673 12621 -2621
rect 12673 -2673 12685 -2621
rect 12737 -2673 12820 -2621
rect 2020 -2680 12820 -2673
rect 2032 -2684 2110 -2680
rect 3980 -2812 4060 -2790
rect 3980 -2868 3992 -2812
rect 4048 -2868 4060 -2812
rect 3980 -2874 3994 -2868
rect 4046 -2874 4060 -2868
rect 3980 -2886 4060 -2874
rect 3980 -2892 3994 -2886
rect 4046 -2892 4060 -2886
rect 3980 -2948 3992 -2892
rect 4048 -2948 4060 -2892
rect 3980 -2970 4060 -2948
rect 5240 -2812 5320 -2790
rect 5240 -2868 5252 -2812
rect 5308 -2868 5320 -2812
rect 5240 -2874 5254 -2868
rect 5306 -2874 5320 -2868
rect 5240 -2886 5320 -2874
rect 5240 -2892 5254 -2886
rect 5306 -2892 5320 -2886
rect 5240 -2948 5252 -2892
rect 5308 -2948 5320 -2892
rect 5240 -2970 5320 -2948
rect 9040 -2812 9120 -2790
rect 9040 -2868 9052 -2812
rect 9108 -2868 9120 -2812
rect 9040 -2874 9054 -2868
rect 9106 -2874 9120 -2868
rect 9040 -2886 9120 -2874
rect 9040 -2892 9054 -2886
rect 9106 -2892 9120 -2886
rect 9040 -2948 9052 -2892
rect 9108 -2948 9120 -2892
rect 9040 -2970 9120 -2948
rect 11560 -2812 11640 -2790
rect 11560 -2868 11572 -2812
rect 11628 -2868 11640 -2812
rect 11560 -2874 11574 -2868
rect 11626 -2874 11640 -2868
rect 11560 -2886 11640 -2874
rect 11560 -2892 11574 -2886
rect 11626 -2892 11640 -2886
rect 11560 -2948 11572 -2892
rect 11628 -2948 11640 -2892
rect 11560 -2970 11640 -2948
rect 12820 -2812 12900 -2790
rect 12820 -2868 12832 -2812
rect 12888 -2868 12900 -2812
rect 12820 -2874 12834 -2868
rect 12886 -2874 12900 -2868
rect 12820 -2886 12900 -2874
rect 12820 -2892 12834 -2886
rect 12886 -2892 12900 -2886
rect 12820 -2948 12832 -2892
rect 12888 -2948 12900 -2892
rect 12820 -2970 12900 -2948
rect 2020 -3090 2100 -3080
rect 2020 -3106 5229 -3090
rect 5440 -3096 6460 -3080
rect 2020 -3158 2032 -3106
rect 2084 -3108 5229 -3106
rect 2084 -3158 2969 -3108
rect 2020 -3160 2969 -3158
rect 3021 -3160 3033 -3108
rect 3085 -3160 3097 -3108
rect 3149 -3160 3161 -3108
rect 3213 -3160 3225 -3108
rect 3277 -3160 3289 -3108
rect 3341 -3160 3353 -3108
rect 3405 -3160 3417 -3108
rect 3469 -3160 3481 -3108
rect 3533 -3160 3545 -3108
rect 3597 -3160 3609 -3108
rect 3661 -3160 3673 -3108
rect 3725 -3160 3737 -3108
rect 3789 -3160 3801 -3108
rect 3853 -3115 5229 -3108
rect 3853 -3160 4248 -3115
rect 2020 -3167 4248 -3160
rect 4300 -3167 4312 -3115
rect 4364 -3167 4376 -3115
rect 4428 -3167 4440 -3115
rect 4492 -3167 4504 -3115
rect 4556 -3167 4568 -3115
rect 4620 -3167 4632 -3115
rect 4684 -3167 4696 -3115
rect 4748 -3167 4760 -3115
rect 4812 -3167 4824 -3115
rect 4876 -3167 4888 -3115
rect 4940 -3167 4952 -3115
rect 5004 -3167 5016 -3115
rect 5068 -3167 5080 -3115
rect 5132 -3167 5229 -3115
rect 2020 -3180 5229 -3167
rect 5260 -3117 5341 -3100
rect 5260 -3169 5273 -3117
rect 5325 -3120 5341 -3117
rect 5440 -3120 5474 -3096
rect 5325 -3148 5474 -3120
rect 5526 -3148 5538 -3096
rect 5590 -3148 5602 -3096
rect 5654 -3148 5666 -3096
rect 5718 -3148 5730 -3096
rect 5782 -3148 5794 -3096
rect 5846 -3148 5858 -3096
rect 5910 -3148 5922 -3096
rect 5974 -3148 5986 -3096
rect 6038 -3148 6050 -3096
rect 6102 -3148 6114 -3096
rect 6166 -3148 6178 -3096
rect 6230 -3148 6242 -3096
rect 6294 -3148 6306 -3096
rect 6358 -3148 6370 -3096
rect 6422 -3148 6460 -3096
rect 5325 -3169 6460 -3148
rect 5260 -3180 6460 -3169
rect 6700 -3103 8980 -3080
rect 9240 -3093 10240 -3080
rect 6700 -3104 7864 -3103
rect 6700 -3156 6726 -3104
rect 6778 -3156 6790 -3104
rect 6842 -3156 6854 -3104
rect 6906 -3156 6918 -3104
rect 6970 -3156 6982 -3104
rect 7034 -3156 7046 -3104
rect 7098 -3156 7110 -3104
rect 7162 -3156 7174 -3104
rect 7226 -3156 7238 -3104
rect 7290 -3156 7302 -3104
rect 7354 -3156 7366 -3104
rect 7418 -3156 7430 -3104
rect 7482 -3156 7494 -3104
rect 7546 -3156 7558 -3104
rect 7610 -3156 7622 -3104
rect 7674 -3156 7864 -3104
rect 6700 -3159 7864 -3156
rect 7920 -3104 8980 -3103
rect 7920 -3156 7986 -3104
rect 8038 -3156 8050 -3104
rect 8102 -3156 8114 -3104
rect 8166 -3156 8178 -3104
rect 8230 -3156 8242 -3104
rect 8294 -3156 8306 -3104
rect 8358 -3156 8370 -3104
rect 8422 -3156 8434 -3104
rect 8486 -3156 8498 -3104
rect 8550 -3156 8562 -3104
rect 8614 -3156 8626 -3104
rect 8678 -3156 8690 -3104
rect 8742 -3156 8754 -3104
rect 8806 -3156 8818 -3104
rect 8870 -3156 8882 -3104
rect 8934 -3156 8980 -3104
rect 7920 -3159 8980 -3156
rect 6700 -3180 8980 -3159
rect 9040 -3116 9120 -3100
rect 9040 -3168 9055 -3116
rect 9107 -3120 9120 -3116
rect 9240 -3120 9264 -3093
rect 9107 -3145 9264 -3120
rect 9316 -3145 9328 -3093
rect 9380 -3145 9392 -3093
rect 9444 -3145 9456 -3093
rect 9508 -3145 9520 -3093
rect 9572 -3145 9584 -3093
rect 9636 -3145 9648 -3093
rect 9700 -3145 9712 -3093
rect 9764 -3145 9776 -3093
rect 9828 -3145 9840 -3093
rect 9892 -3145 9904 -3093
rect 9956 -3145 9968 -3093
rect 10020 -3145 10032 -3093
rect 10084 -3145 10096 -3093
rect 10148 -3145 10160 -3093
rect 10212 -3145 10240 -3093
rect 9107 -3168 10240 -3145
rect 9040 -3180 10240 -3168
rect 10311 -3104 10368 -3089
rect 10311 -3134 10313 -3104
rect 10365 -3134 10368 -3104
rect 5269 -3183 5329 -3180
rect 9050 -3182 9113 -3180
rect 10367 -3190 10368 -3134
rect 10500 -3103 13630 -3090
rect 10500 -3108 11812 -3103
rect 10500 -3160 10553 -3108
rect 10605 -3160 10617 -3108
rect 10669 -3160 10681 -3108
rect 10733 -3160 10745 -3108
rect 10797 -3160 10809 -3108
rect 10861 -3160 10873 -3108
rect 10925 -3160 10937 -3108
rect 10989 -3160 11001 -3108
rect 11053 -3160 11065 -3108
rect 11117 -3160 11129 -3108
rect 11181 -3160 11193 -3108
rect 11245 -3160 11257 -3108
rect 11309 -3160 11321 -3108
rect 11373 -3160 11385 -3108
rect 11437 -3155 11812 -3108
rect 11864 -3155 11876 -3103
rect 11928 -3155 11940 -3103
rect 11992 -3155 12004 -3103
rect 12056 -3155 12068 -3103
rect 12120 -3155 12132 -3103
rect 12184 -3155 12196 -3103
rect 12248 -3155 12260 -3103
rect 12312 -3155 12324 -3103
rect 12376 -3155 12388 -3103
rect 12440 -3155 12452 -3103
rect 12504 -3155 12516 -3103
rect 12568 -3155 12580 -3103
rect 12632 -3155 12644 -3103
rect 12696 -3112 13630 -3103
rect 12696 -3155 13564 -3112
rect 11437 -3160 13564 -3155
rect 10500 -3164 13564 -3160
rect 13616 -3164 13630 -3112
rect 10500 -3180 13630 -3164
rect 10311 -3220 10313 -3190
rect 10365 -3220 10368 -3190
rect 10311 -3234 10368 -3220
rect 2020 -3866 9450 -3850
rect 2020 -3882 2776 -3866
rect 2020 -3938 2052 -3882
rect 2108 -3892 2776 -3882
rect 2108 -3897 2419 -3892
rect 2108 -3938 2294 -3897
rect 2020 -3949 2294 -3938
rect 2346 -3944 2419 -3897
rect 2471 -3918 2776 -3892
rect 2828 -3904 9450 -3866
rect 2828 -3918 9384 -3904
rect 2471 -3930 9384 -3918
rect 2471 -3944 2776 -3930
rect 2346 -3949 2776 -3944
rect 2020 -3956 2776 -3949
rect 2020 -3961 2419 -3956
rect 2020 -3962 2294 -3961
rect 2020 -4018 2052 -3962
rect 2108 -4013 2294 -3962
rect 2346 -4008 2419 -3961
rect 2471 -3982 2776 -3956
rect 2828 -3956 9384 -3930
rect 9436 -3956 9450 -3904
rect 2828 -3982 9450 -3956
rect 2471 -3994 9450 -3982
rect 2471 -4008 2776 -3994
rect 2346 -4013 2776 -4008
rect 2108 -4018 2776 -4013
rect 2020 -4046 2776 -4018
rect 2828 -4046 9384 -3994
rect 9436 -4046 9450 -3994
rect 2020 -4060 9450 -4046
rect 2870 -4103 10380 -4090
rect 2870 -4104 10311 -4103
rect 2870 -4156 2879 -4104
rect 2931 -4156 9494 -4104
rect 9546 -4156 9574 -4104
rect 9626 -4156 10311 -4104
rect 2870 -4159 10311 -4156
rect 10367 -4159 10380 -4103
rect 2870 -4170 10380 -4159
rect 10311 -4172 10368 -4170
rect 2150 -4213 13960 -4200
rect 2150 -4265 2163 -4213
rect 2215 -4214 13960 -4213
rect 2215 -4265 13566 -4214
rect 2150 -4266 13566 -4265
rect 13618 -4266 13960 -4214
rect 2150 -4280 13960 -4266
rect 1780 -4323 13960 -4310
rect 1780 -4375 1794 -4323
rect 1846 -4328 13960 -4323
rect 1846 -4375 13674 -4328
rect 1780 -4380 13674 -4375
rect 13726 -4380 13960 -4328
rect 1780 -4390 13960 -4380
rect 1670 -4432 13960 -4420
rect 1670 -4433 13782 -4432
rect 1670 -4485 1681 -4433
rect 1733 -4484 13782 -4433
rect 13834 -4484 13960 -4432
rect 1733 -4485 13960 -4484
rect 1670 -4500 13960 -4485
rect 2020 -4546 13960 -4530
rect 2020 -4598 2034 -4546
rect 2086 -4598 13894 -4546
rect 13946 -4598 13960 -4546
rect 2020 -4610 13960 -4598
rect 2980 -4652 7940 -4640
rect 2980 -4655 7852 -4652
rect 2980 -4707 2995 -4655
rect 3047 -4707 7852 -4655
rect 2980 -4708 7852 -4707
rect 7908 -4708 7940 -4652
rect 2980 -4720 7940 -4708
rect 6461 -4721 6559 -4720
rect 1890 -4772 2070 -4740
rect 7802 -4759 8705 -4757
rect 7802 -4760 8801 -4759
rect 1890 -4828 1912 -4772
rect 1968 -4828 2070 -4772
rect 1890 -4836 2070 -4828
rect 1890 -4862 1914 -4836
rect 1966 -4862 2070 -4836
rect 1890 -4918 1912 -4862
rect 1968 -4918 2070 -4862
rect 1890 -4940 2070 -4918
rect 2760 -4782 8801 -4760
rect 2760 -4787 8622 -4782
rect 2760 -4792 6652 -4787
rect 2760 -4848 4912 -4792
rect 4968 -4848 6072 -4792
rect 6128 -4848 6152 -4792
rect 6208 -4843 6652 -4792
rect 6708 -4843 7472 -4787
rect 7528 -4838 8622 -4787
rect 8678 -4838 8801 -4782
rect 7528 -4843 8801 -4838
rect 6208 -4848 8801 -4843
rect 2760 -4869 8801 -4848
rect 2760 -4870 6250 -4869
rect 7350 -4870 7470 -4869
rect 2760 -4950 2850 -4870
rect 6030 -4880 6250 -4870
rect 2100 -4954 2850 -4950
rect 2100 -5006 2149 -4954
rect 2201 -5006 2289 -4954
rect 2341 -5006 2419 -4954
rect 2471 -5006 2850 -4954
rect 2100 -5030 2850 -5006
rect 4804 -5510 4863 -5506
rect 6056 -5509 6115 -5506
rect 6056 -5510 6121 -5509
rect 7299 -5510 7358 -5505
rect 8534 -5510 8605 -5505
rect 2980 -5521 8610 -5510
rect 2980 -5522 7302 -5521
rect 2980 -5526 4807 -5522
rect 2980 -5578 2996 -5526
rect 3048 -5547 4807 -5526
rect 3048 -5578 4126 -5547
rect 2980 -5590 4126 -5578
rect 2993 -5593 3052 -5590
rect 4102 -5599 4126 -5590
rect 4178 -5599 4190 -5547
rect 4242 -5599 4254 -5547
rect 4306 -5599 4318 -5547
rect 4370 -5599 4382 -5547
rect 4434 -5574 4807 -5547
rect 4859 -5543 6059 -5522
rect 4859 -5574 5413 -5543
rect 4434 -5590 5413 -5574
rect 4434 -5599 4458 -5590
rect 4102 -5617 4458 -5599
rect 5389 -5595 5413 -5590
rect 5465 -5595 5477 -5543
rect 5529 -5595 5541 -5543
rect 5593 -5595 5605 -5543
rect 5657 -5595 5669 -5543
rect 5721 -5574 6059 -5543
rect 6111 -5545 7302 -5522
rect 6111 -5574 6693 -5545
rect 5721 -5590 6693 -5574
rect 5721 -5595 5745 -5590
rect 5389 -5613 5745 -5595
rect 6669 -5597 6693 -5590
rect 6745 -5597 6757 -5545
rect 6809 -5597 6821 -5545
rect 6873 -5597 6885 -5545
rect 6937 -5597 6949 -5545
rect 7001 -5573 7302 -5545
rect 7354 -5522 8610 -5521
rect 7354 -5547 8543 -5522
rect 7354 -5573 7928 -5547
rect 7001 -5590 7928 -5573
rect 7001 -5597 7025 -5590
rect 6669 -5615 7025 -5597
rect 7904 -5599 7928 -5590
rect 7980 -5599 7992 -5547
rect 8044 -5599 8056 -5547
rect 8108 -5599 8120 -5547
rect 8172 -5599 8184 -5547
rect 8236 -5574 8543 -5547
rect 8595 -5574 8610 -5522
rect 8236 -5590 8610 -5574
rect 8236 -5599 8260 -5590
rect 7904 -5617 8260 -5599
rect 3750 -6059 9670 -6050
rect 3750 -6062 3802 -6059
rect 3854 -6062 3866 -6059
rect 3750 -6118 3762 -6062
rect 3918 -6111 3930 -6059
rect 3982 -6111 3994 -6059
rect 4046 -6111 4058 -6059
rect 4110 -6111 4122 -6059
rect 4174 -6111 4186 -6059
rect 4238 -6111 4250 -6059
rect 4302 -6111 4314 -6059
rect 4366 -6111 4378 -6059
rect 4430 -6111 4442 -6059
rect 4494 -6111 4506 -6059
rect 4558 -6111 4570 -6059
rect 4622 -6111 4634 -6059
rect 4686 -6061 9670 -6059
rect 4686 -6063 6275 -6061
rect 4686 -6111 5031 -6063
rect 3818 -6118 3852 -6111
rect 3908 -6115 5031 -6111
rect 5083 -6115 5095 -6063
rect 5147 -6115 5159 -6063
rect 5211 -6115 5223 -6063
rect 5275 -6115 5287 -6063
rect 5339 -6115 5351 -6063
rect 5403 -6115 5415 -6063
rect 5467 -6115 5479 -6063
rect 5531 -6115 5543 -6063
rect 5595 -6115 5607 -6063
rect 5659 -6115 5671 -6063
rect 5723 -6115 5735 -6063
rect 5787 -6115 5799 -6063
rect 5851 -6115 5863 -6063
rect 5915 -6115 5927 -6063
rect 5979 -6113 6275 -6063
rect 6327 -6113 6339 -6061
rect 6391 -6113 6403 -6061
rect 6455 -6113 6467 -6061
rect 6519 -6113 6531 -6061
rect 6583 -6113 6595 -6061
rect 6647 -6113 6659 -6061
rect 6711 -6113 6723 -6061
rect 6775 -6113 6787 -6061
rect 6839 -6113 6851 -6061
rect 6903 -6113 6915 -6061
rect 6967 -6113 6979 -6061
rect 7031 -6113 7043 -6061
rect 7095 -6113 7107 -6061
rect 7159 -6113 7171 -6061
rect 7223 -6064 9670 -6061
rect 7223 -6066 9604 -6064
rect 7223 -6113 7513 -6066
rect 5979 -6115 7513 -6113
rect 3908 -6118 7513 -6115
rect 7565 -6118 7577 -6066
rect 7629 -6118 7641 -6066
rect 7693 -6118 7705 -6066
rect 7757 -6118 7769 -6066
rect 7821 -6118 7833 -6066
rect 7885 -6118 7897 -6066
rect 7949 -6118 7961 -6066
rect 8013 -6118 8025 -6066
rect 8077 -6118 8089 -6066
rect 8141 -6118 8153 -6066
rect 8205 -6118 8217 -6066
rect 8269 -6118 8281 -6066
rect 8333 -6118 8345 -6066
rect 8397 -6118 8409 -6066
rect 8461 -6116 9604 -6066
rect 9656 -6116 9670 -6064
rect 8461 -6118 9670 -6116
rect 3750 -6130 9670 -6118
rect 2760 -6216 2870 -6210
rect 3060 -6216 3770 -6210
rect 2760 -6234 4674 -6216
rect 2760 -6286 2774 -6234
rect 2826 -6250 4674 -6234
rect 2826 -6286 3793 -6250
rect 2760 -6302 3793 -6286
rect 3845 -6302 3857 -6250
rect 3909 -6302 3921 -6250
rect 3973 -6302 3985 -6250
rect 4037 -6302 4049 -6250
rect 4101 -6302 4113 -6250
rect 4165 -6302 4177 -6250
rect 4229 -6302 4241 -6250
rect 4293 -6302 4305 -6250
rect 4357 -6302 4369 -6250
rect 4421 -6302 4674 -6250
rect 5110 -6225 5895 -6210
rect 8670 -6214 9560 -6210
rect 5110 -6281 5114 -6225
rect 5170 -6227 5194 -6225
rect 5250 -6227 5274 -6225
rect 5330 -6227 5354 -6225
rect 5410 -6227 5434 -6225
rect 5490 -6227 5514 -6225
rect 5570 -6227 5594 -6225
rect 5650 -6227 5674 -6225
rect 5730 -6227 5754 -6225
rect 5810 -6227 5834 -6225
rect 5176 -6279 5188 -6227
rect 5250 -6279 5252 -6227
rect 5432 -6279 5434 -6227
rect 5496 -6279 5508 -6227
rect 5570 -6279 5572 -6227
rect 5752 -6279 5754 -6227
rect 5816 -6279 5828 -6227
rect 5170 -6281 5194 -6279
rect 5250 -6281 5274 -6279
rect 5330 -6281 5354 -6279
rect 5410 -6281 5434 -6279
rect 5490 -6281 5514 -6279
rect 5570 -6281 5594 -6279
rect 5650 -6281 5674 -6279
rect 5730 -6281 5754 -6279
rect 5810 -6281 5834 -6279
rect 5890 -6281 5895 -6225
rect 5110 -6296 5895 -6281
rect 7493 -6233 9560 -6214
rect 7493 -6285 7704 -6233
rect 7756 -6285 7768 -6233
rect 7820 -6285 7832 -6233
rect 7884 -6285 7896 -6233
rect 7948 -6285 7960 -6233
rect 8012 -6285 8024 -6233
rect 8076 -6285 8088 -6233
rect 8140 -6285 8152 -6233
rect 8204 -6285 8216 -6233
rect 8268 -6285 8280 -6233
rect 8332 -6234 9560 -6233
rect 8332 -6285 9494 -6234
rect 7493 -6286 9494 -6285
rect 9546 -6286 9560 -6234
rect 2760 -6310 4674 -6302
rect 7493 -6310 9560 -6286
rect 3771 -6317 4443 -6310
rect 7493 -6312 8710 -6310
rect 9510 -6312 9560 -6310
rect 6104 -6370 6175 -6357
rect 6104 -6376 6113 -6370
rect 6165 -6376 6175 -6370
rect 4800 -6458 4869 -6428
rect 4800 -6514 4806 -6458
rect 4862 -6514 4869 -6458
rect 4800 -6520 4808 -6514
rect 4860 -6520 4869 -6514
rect 4800 -6532 4869 -6520
rect 4800 -6538 4808 -6532
rect 4860 -6538 4869 -6532
rect 4800 -6594 4806 -6538
rect 4862 -6594 4869 -6538
rect 4800 -6623 4869 -6594
rect 6104 -6432 6111 -6376
rect 6167 -6432 6175 -6376
rect 6104 -6434 6175 -6432
rect 6104 -6456 6113 -6434
rect 6165 -6456 6175 -6434
rect 6104 -6512 6111 -6456
rect 6167 -6512 6175 -6456
rect 6104 -6536 6113 -6512
rect 6165 -6536 6175 -6512
rect 6104 -6592 6111 -6536
rect 6167 -6592 6175 -6536
rect 6104 -6614 6113 -6592
rect 6165 -6614 6175 -6592
rect 6104 -6616 6175 -6614
rect 6104 -6672 6111 -6616
rect 6167 -6672 6175 -6616
rect 6104 -6678 6113 -6672
rect 6165 -6678 6175 -6672
rect 6104 -6690 6175 -6678
rect 7362 -6365 7433 -6352
rect 7362 -6371 7371 -6365
rect 7423 -6371 7433 -6365
rect 7362 -6427 7369 -6371
rect 7425 -6427 7433 -6371
rect 7362 -6429 7433 -6427
rect 7362 -6451 7371 -6429
rect 7423 -6451 7433 -6429
rect 7362 -6507 7369 -6451
rect 7425 -6507 7433 -6451
rect 7362 -6531 7371 -6507
rect 7423 -6531 7433 -6507
rect 7362 -6587 7369 -6531
rect 7425 -6587 7433 -6531
rect 7362 -6609 7371 -6587
rect 7423 -6609 7433 -6587
rect 7362 -6611 7433 -6609
rect 7362 -6667 7369 -6611
rect 7425 -6667 7433 -6611
rect 7362 -6673 7371 -6667
rect 7423 -6673 7433 -6667
rect 7362 -6685 7433 -6673
rect 2670 -6742 8510 -6730
rect 2670 -6746 3781 -6742
rect 2670 -6798 2681 -6746
rect 2733 -6794 3781 -6746
rect 3833 -6794 3845 -6742
rect 3897 -6794 3909 -6742
rect 3961 -6794 3973 -6742
rect 4025 -6794 4037 -6742
rect 4089 -6794 4101 -6742
rect 4153 -6794 4165 -6742
rect 4217 -6794 4229 -6742
rect 4281 -6794 4293 -6742
rect 4345 -6794 4357 -6742
rect 4409 -6794 4421 -6742
rect 4473 -6794 4485 -6742
rect 4537 -6794 4549 -6742
rect 4601 -6794 4613 -6742
rect 4665 -6794 4677 -6742
rect 4729 -6745 7513 -6742
rect 4729 -6748 6281 -6745
rect 4729 -6794 5024 -6748
rect 2733 -6798 5024 -6794
rect 2670 -6800 5024 -6798
rect 5076 -6800 5088 -6748
rect 5140 -6800 5152 -6748
rect 5204 -6800 5216 -6748
rect 5268 -6800 5280 -6748
rect 5332 -6800 5344 -6748
rect 5396 -6800 5408 -6748
rect 5460 -6800 5472 -6748
rect 5524 -6800 5536 -6748
rect 5588 -6800 5600 -6748
rect 5652 -6800 5664 -6748
rect 5716 -6800 5728 -6748
rect 5780 -6800 5792 -6748
rect 5844 -6800 5856 -6748
rect 5908 -6800 5920 -6748
rect 5972 -6797 6281 -6748
rect 6333 -6797 6345 -6745
rect 6397 -6797 6409 -6745
rect 6461 -6797 6473 -6745
rect 6525 -6797 6537 -6745
rect 6589 -6797 6601 -6745
rect 6653 -6797 6665 -6745
rect 6717 -6797 6729 -6745
rect 6781 -6797 6793 -6745
rect 6845 -6797 6857 -6745
rect 6909 -6797 6921 -6745
rect 6973 -6797 6985 -6745
rect 7037 -6797 7049 -6745
rect 7101 -6797 7113 -6745
rect 7165 -6797 7177 -6745
rect 7229 -6794 7513 -6745
rect 7565 -6794 7577 -6742
rect 7629 -6794 7641 -6742
rect 7693 -6794 7705 -6742
rect 7757 -6794 7769 -6742
rect 7821 -6794 7833 -6742
rect 7885 -6794 7897 -6742
rect 7949 -6794 7961 -6742
rect 8013 -6794 8025 -6742
rect 8077 -6794 8089 -6742
rect 8141 -6794 8153 -6742
rect 8205 -6794 8217 -6742
rect 8269 -6794 8281 -6742
rect 8333 -6794 8345 -6742
rect 8397 -6794 8409 -6742
rect 8461 -6794 8510 -6742
rect 7229 -6797 8510 -6794
rect 5972 -6800 8510 -6797
rect 2670 -6810 8510 -6800
rect 6390 -6909 7175 -6894
rect 2870 -6924 4750 -6910
rect 2870 -6976 2884 -6924
rect 2936 -6926 4750 -6924
rect 2936 -6976 3792 -6926
rect 2870 -6978 3792 -6976
rect 3844 -6978 3856 -6926
rect 3908 -6978 3920 -6926
rect 3972 -6978 3984 -6926
rect 4036 -6978 4048 -6926
rect 4100 -6978 4112 -6926
rect 4164 -6978 4176 -6926
rect 4228 -6978 4240 -6926
rect 4292 -6978 4304 -6926
rect 4356 -6978 4368 -6926
rect 4420 -6978 4750 -6926
rect 2870 -6990 4750 -6978
rect 6390 -6965 6394 -6909
rect 6450 -6911 6474 -6909
rect 6530 -6911 6554 -6909
rect 6610 -6911 6634 -6909
rect 6690 -6911 6714 -6909
rect 6770 -6911 6794 -6909
rect 6850 -6911 6874 -6909
rect 6930 -6911 6954 -6909
rect 7010 -6911 7034 -6909
rect 7090 -6911 7114 -6909
rect 6456 -6963 6468 -6911
rect 6530 -6963 6532 -6911
rect 6712 -6963 6714 -6911
rect 6776 -6963 6788 -6911
rect 6850 -6963 6852 -6911
rect 7032 -6963 7034 -6911
rect 7096 -6963 7108 -6911
rect 6450 -6965 6474 -6963
rect 6530 -6965 6554 -6963
rect 6610 -6965 6634 -6963
rect 6690 -6965 6714 -6963
rect 6770 -6965 6794 -6963
rect 6850 -6965 6874 -6963
rect 6930 -6965 6954 -6963
rect 7010 -6965 7034 -6963
rect 7090 -6965 7114 -6963
rect 7170 -6965 7175 -6909
rect 7637 -6910 8309 -6909
rect 6390 -6980 7175 -6965
rect 7493 -6924 9450 -6910
rect 7493 -6925 9385 -6924
rect 7493 -6977 7659 -6925
rect 7711 -6977 7723 -6925
rect 7775 -6977 7787 -6925
rect 7839 -6977 7851 -6925
rect 7903 -6977 7915 -6925
rect 7967 -6977 7979 -6925
rect 8031 -6977 8043 -6925
rect 8095 -6977 8107 -6925
rect 8159 -6977 8171 -6925
rect 8223 -6977 8235 -6925
rect 8287 -6976 9385 -6925
rect 9437 -6976 9450 -6924
rect 8287 -6977 9450 -6976
rect 7493 -6986 9450 -6977
rect 3770 -6993 4442 -6990
rect 7637 -6992 8309 -6986
rect 8610 -6990 9450 -6986
rect 8610 -7032 8690 -7020
rect 8610 -7088 8622 -7032
rect 8678 -7088 8690 -7032
rect 8610 -7110 8624 -7088
rect 8676 -7110 8690 -7088
rect 8610 -7112 8690 -7110
rect 8610 -7168 8622 -7112
rect 8678 -7168 8690 -7112
rect 8610 -7174 8624 -7168
rect 8676 -7174 8690 -7168
rect 8610 -7186 8690 -7174
rect 8610 -7192 8624 -7186
rect 8676 -7192 8690 -7186
rect 8610 -7248 8622 -7192
rect 8678 -7248 8690 -7192
rect 8610 -7250 8690 -7248
rect 8610 -7272 8624 -7250
rect 8676 -7272 8690 -7250
rect 8610 -7328 8622 -7272
rect 8678 -7328 8690 -7272
rect 8610 -7340 8690 -7328
rect 2670 -7421 8510 -7410
rect 2670 -7424 3775 -7421
rect 2670 -7476 2689 -7424
rect 2741 -7473 3775 -7424
rect 3827 -7473 3839 -7421
rect 3891 -7473 3903 -7421
rect 3955 -7473 3967 -7421
rect 4019 -7473 4031 -7421
rect 4083 -7473 4095 -7421
rect 4147 -7473 4159 -7421
rect 4211 -7473 4223 -7421
rect 4275 -7473 4287 -7421
rect 4339 -7473 4351 -7421
rect 4403 -7473 4415 -7421
rect 4467 -7473 4479 -7421
rect 4531 -7473 4543 -7421
rect 4595 -7473 4607 -7421
rect 4659 -7473 4671 -7421
rect 4723 -7473 5014 -7421
rect 5066 -7473 5078 -7421
rect 5130 -7473 5142 -7421
rect 5194 -7473 5206 -7421
rect 5258 -7473 5270 -7421
rect 5322 -7473 5334 -7421
rect 5386 -7473 5398 -7421
rect 5450 -7473 5462 -7421
rect 5514 -7473 5526 -7421
rect 5578 -7473 5590 -7421
rect 5642 -7473 5654 -7421
rect 5706 -7473 5718 -7421
rect 5770 -7473 5782 -7421
rect 5834 -7473 5846 -7421
rect 5898 -7473 5910 -7421
rect 5962 -7422 8510 -7421
rect 5962 -7425 7516 -7422
rect 5962 -7473 6256 -7425
rect 2741 -7476 6256 -7473
rect 2670 -7477 6256 -7476
rect 6308 -7477 6320 -7425
rect 6372 -7477 6384 -7425
rect 6436 -7477 6448 -7425
rect 6500 -7477 6512 -7425
rect 6564 -7477 6576 -7425
rect 6628 -7477 6640 -7425
rect 6692 -7477 6704 -7425
rect 6756 -7477 6768 -7425
rect 6820 -7477 6832 -7425
rect 6884 -7477 6896 -7425
rect 6948 -7477 6960 -7425
rect 7012 -7477 7024 -7425
rect 7076 -7477 7088 -7425
rect 7140 -7477 7152 -7425
rect 7204 -7474 7516 -7425
rect 7568 -7474 7580 -7422
rect 7632 -7474 7644 -7422
rect 7696 -7474 7708 -7422
rect 7760 -7474 7772 -7422
rect 7824 -7474 7836 -7422
rect 7888 -7474 7900 -7422
rect 7952 -7474 7964 -7422
rect 8016 -7474 8028 -7422
rect 8080 -7474 8092 -7422
rect 8144 -7474 8156 -7422
rect 8208 -7474 8220 -7422
rect 8272 -7474 8284 -7422
rect 8336 -7474 8348 -7422
rect 8400 -7474 8412 -7422
rect 8464 -7474 8510 -7422
rect 7204 -7477 8510 -7474
rect 2670 -7490 8510 -7477
rect 2980 -7596 8610 -7590
rect 2980 -7604 4112 -7596
rect 2980 -7656 2994 -7604
rect 3046 -7648 4112 -7604
rect 4164 -7648 4176 -7596
rect 4228 -7648 4240 -7596
rect 4292 -7648 4304 -7596
rect 4356 -7604 5340 -7596
rect 4356 -7648 4802 -7604
rect 3046 -7656 4802 -7648
rect 4854 -7648 5340 -7604
rect 5392 -7648 5404 -7596
rect 5456 -7648 5468 -7596
rect 5520 -7648 5532 -7596
rect 5584 -7597 8610 -7596
rect 5584 -7601 7905 -7597
rect 5584 -7605 6637 -7601
rect 5584 -7648 6041 -7605
rect 4854 -7656 6041 -7648
rect 2980 -7657 6041 -7656
rect 6093 -7653 6637 -7605
rect 6689 -7653 6701 -7601
rect 6753 -7653 6765 -7601
rect 6817 -7653 6829 -7601
rect 6881 -7611 7905 -7601
rect 6881 -7653 7281 -7611
rect 6093 -7657 7281 -7653
rect 2980 -7663 7281 -7657
rect 7333 -7649 7905 -7611
rect 7957 -7649 7969 -7597
rect 8021 -7649 8033 -7597
rect 8085 -7649 8097 -7597
rect 8149 -7605 8610 -7597
rect 8149 -7649 8545 -7605
rect 7333 -7657 8545 -7649
rect 8597 -7657 8610 -7605
rect 7333 -7663 8610 -7657
rect 2980 -7670 8610 -7663
rect 3750 -8098 9670 -8090
rect 3750 -8104 6259 -8098
rect 3750 -8156 3778 -8104
rect 3830 -8156 3842 -8104
rect 3894 -8156 3906 -8104
rect 3958 -8156 3970 -8104
rect 4022 -8156 4034 -8104
rect 4086 -8156 4098 -8104
rect 4150 -8156 4162 -8104
rect 4214 -8156 4226 -8104
rect 4278 -8156 4290 -8104
rect 4342 -8156 4354 -8104
rect 4406 -8156 4418 -8104
rect 4470 -8156 4482 -8104
rect 4534 -8156 4546 -8104
rect 4598 -8156 4610 -8104
rect 4662 -8156 4674 -8104
rect 4726 -8156 5020 -8104
rect 5072 -8156 5084 -8104
rect 5136 -8156 5148 -8104
rect 5200 -8156 5212 -8104
rect 5264 -8156 5276 -8104
rect 5328 -8156 5340 -8104
rect 5392 -8156 5404 -8104
rect 5456 -8156 5468 -8104
rect 5520 -8156 5532 -8104
rect 5584 -8156 5596 -8104
rect 5648 -8156 5660 -8104
rect 5712 -8156 5724 -8104
rect 5776 -8156 5788 -8104
rect 5840 -8156 5852 -8104
rect 5904 -8156 5916 -8104
rect 5968 -8150 6259 -8104
rect 6311 -8150 6323 -8098
rect 6375 -8150 6387 -8098
rect 6439 -8150 6451 -8098
rect 6503 -8150 6515 -8098
rect 6567 -8150 6579 -8098
rect 6631 -8150 6643 -8098
rect 6695 -8150 6707 -8098
rect 6759 -8150 6771 -8098
rect 6823 -8150 6835 -8098
rect 6887 -8150 6899 -8098
rect 6951 -8150 6963 -8098
rect 7015 -8150 7027 -8098
rect 7079 -8150 7091 -8098
rect 7143 -8150 7155 -8098
rect 7207 -8103 9670 -8098
rect 7207 -8150 7521 -8103
rect 5968 -8155 7521 -8150
rect 7573 -8155 7585 -8103
rect 7637 -8155 7649 -8103
rect 7701 -8155 7713 -8103
rect 7765 -8155 7777 -8103
rect 7829 -8155 7841 -8103
rect 7893 -8155 7905 -8103
rect 7957 -8155 7969 -8103
rect 8021 -8155 8033 -8103
rect 8085 -8155 8097 -8103
rect 8149 -8155 8161 -8103
rect 8213 -8155 8225 -8103
rect 8277 -8155 8289 -8103
rect 8341 -8155 8353 -8103
rect 8405 -8155 8417 -8103
rect 8469 -8104 9670 -8103
rect 8469 -8155 9604 -8104
rect 5968 -8156 9604 -8155
rect 9656 -8156 9670 -8104
rect 3750 -8170 9670 -8156
<< via2 >>
rect 6562 72 6618 128
rect 10352 72 10408 128
rect 7652 -388 7708 -332
rect 7652 -468 7708 -412
rect 3992 -762 4048 -752
rect 3992 -808 3994 -762
rect 3994 -808 4046 -762
rect 4046 -808 4048 -762
rect 3992 -878 3994 -832
rect 3994 -878 4046 -832
rect 4046 -878 4048 -832
rect 3992 -888 4048 -878
rect 5252 -762 5308 -752
rect 5252 -808 5254 -762
rect 5254 -808 5306 -762
rect 5306 -808 5308 -762
rect 5252 -878 5254 -832
rect 5254 -878 5306 -832
rect 5306 -878 5308 -832
rect 5252 -888 5308 -878
rect 6562 -708 6618 -682
rect 6562 -738 6564 -708
rect 6564 -738 6616 -708
rect 6616 -738 6618 -708
rect 6562 -772 6618 -762
rect 6562 -818 6564 -772
rect 6564 -818 6616 -772
rect 6616 -818 6618 -772
rect 6562 -888 6564 -842
rect 6564 -888 6616 -842
rect 6616 -888 6618 -842
rect 6562 -898 6618 -888
rect 7772 -762 7828 -752
rect 7772 -808 7774 -762
rect 7774 -808 7826 -762
rect 7826 -808 7828 -762
rect 7772 -878 7774 -832
rect 7774 -878 7826 -832
rect 7826 -878 7828 -832
rect 7772 -888 7828 -878
rect 9032 -762 9088 -752
rect 9032 -808 9034 -762
rect 9034 -808 9086 -762
rect 9086 -808 9088 -762
rect 9032 -878 9034 -832
rect 9034 -878 9086 -832
rect 9086 -878 9088 -832
rect 9032 -888 9088 -878
rect 10354 -776 10356 -738
rect 10356 -776 10408 -738
rect 10408 -776 10410 -738
rect 10354 -788 10410 -776
rect 10354 -794 10356 -788
rect 10356 -794 10408 -788
rect 10408 -794 10410 -788
rect 10354 -840 10356 -818
rect 10356 -840 10408 -818
rect 10408 -840 10410 -818
rect 10354 -852 10410 -840
rect 10354 -874 10356 -852
rect 10356 -874 10408 -852
rect 10408 -874 10410 -852
rect 6562 -952 6564 -922
rect 6564 -952 6616 -922
rect 6616 -952 6618 -922
rect 6562 -978 6618 -952
rect 10354 -904 10356 -898
rect 10356 -904 10408 -898
rect 10408 -904 10410 -898
rect 10354 -916 10410 -904
rect 10354 -954 10356 -916
rect 10356 -954 10408 -916
rect 10408 -954 10410 -916
rect 11572 -762 11628 -752
rect 11572 -808 11574 -762
rect 11574 -808 11626 -762
rect 11626 -808 11628 -762
rect 11572 -878 11574 -832
rect 11574 -878 11626 -832
rect 11626 -878 11628 -832
rect 11572 -888 11628 -878
rect 12832 -762 12888 -752
rect 12832 -808 12834 -762
rect 12834 -808 12886 -762
rect 12886 -808 12888 -762
rect 12832 -878 12834 -832
rect 12834 -878 12886 -832
rect 12886 -878 12888 -832
rect 12832 -888 12888 -878
rect 7853 -1115 7909 -1059
rect 3992 -1462 4048 -1452
rect 3992 -1508 3994 -1462
rect 3994 -1508 4046 -1462
rect 4046 -1508 4048 -1462
rect 3992 -1578 3994 -1532
rect 3994 -1578 4046 -1532
rect 4046 -1578 4048 -1532
rect 3992 -1588 4048 -1578
rect 5272 -1462 5328 -1452
rect 5272 -1508 5274 -1462
rect 5274 -1508 5326 -1462
rect 5326 -1508 5328 -1462
rect 5272 -1578 5274 -1532
rect 5274 -1578 5326 -1532
rect 5326 -1578 5328 -1532
rect 5272 -1588 5328 -1578
rect 9052 -1462 9108 -1452
rect 9052 -1508 9054 -1462
rect 9054 -1508 9106 -1462
rect 9106 -1508 9108 -1462
rect 9052 -1578 9054 -1532
rect 9054 -1578 9106 -1532
rect 9106 -1578 9108 -1532
rect 9052 -1588 9108 -1578
rect 11572 -1462 11628 -1452
rect 11572 -1508 11574 -1462
rect 11574 -1508 11626 -1462
rect 11626 -1508 11628 -1462
rect 11572 -1578 11574 -1532
rect 11574 -1578 11626 -1532
rect 11626 -1578 11628 -1532
rect 11572 -1588 11628 -1578
rect 12832 -1462 12888 -1452
rect 12832 -1508 12834 -1462
rect 12834 -1508 12886 -1462
rect 12886 -1508 12888 -1462
rect 12832 -1578 12834 -1532
rect 12834 -1578 12886 -1532
rect 12886 -1578 12888 -1532
rect 12832 -1588 12888 -1578
rect 6649 -1809 6705 -1753
rect 3992 -2162 4048 -2152
rect 3992 -2208 3994 -2162
rect 3994 -2208 4046 -2162
rect 4046 -2208 4048 -2162
rect 3992 -2278 3994 -2232
rect 3994 -2278 4046 -2232
rect 4046 -2278 4048 -2232
rect 3992 -2288 4048 -2278
rect 5252 -2162 5308 -2152
rect 5252 -2208 5254 -2162
rect 5254 -2208 5306 -2162
rect 5306 -2208 5308 -2162
rect 5252 -2278 5254 -2232
rect 5254 -2278 5306 -2232
rect 5306 -2278 5308 -2232
rect 5252 -2288 5308 -2278
rect 9052 -2162 9108 -2152
rect 9052 -2208 9054 -2162
rect 9054 -2208 9106 -2162
rect 9106 -2208 9108 -2162
rect 9052 -2278 9054 -2232
rect 9054 -2278 9106 -2232
rect 9106 -2278 9108 -2232
rect 9052 -2288 9108 -2278
rect 11572 -2162 11628 -2152
rect 11572 -2208 11574 -2162
rect 11574 -2208 11626 -2162
rect 11626 -2208 11628 -2162
rect 11572 -2278 11574 -2232
rect 11574 -2278 11626 -2232
rect 11626 -2278 11628 -2232
rect 11572 -2288 11628 -2278
rect 12832 -2162 12888 -2152
rect 12832 -2208 12834 -2162
rect 12834 -2208 12886 -2162
rect 12886 -2208 12888 -2162
rect 12832 -2278 12834 -2232
rect 12834 -2278 12886 -2232
rect 12886 -2278 12888 -2232
rect 12832 -2288 12888 -2278
rect 6651 -2490 6707 -2434
rect 3992 -2822 4048 -2812
rect 3992 -2868 3994 -2822
rect 3994 -2868 4046 -2822
rect 4046 -2868 4048 -2822
rect 3992 -2938 3994 -2892
rect 3994 -2938 4046 -2892
rect 4046 -2938 4048 -2892
rect 3992 -2948 4048 -2938
rect 5252 -2822 5308 -2812
rect 5252 -2868 5254 -2822
rect 5254 -2868 5306 -2822
rect 5306 -2868 5308 -2822
rect 5252 -2938 5254 -2892
rect 5254 -2938 5306 -2892
rect 5306 -2938 5308 -2892
rect 5252 -2948 5308 -2938
rect 9052 -2822 9108 -2812
rect 9052 -2868 9054 -2822
rect 9054 -2868 9106 -2822
rect 9106 -2868 9108 -2822
rect 9052 -2938 9054 -2892
rect 9054 -2938 9106 -2892
rect 9106 -2938 9108 -2892
rect 9052 -2948 9108 -2938
rect 11572 -2822 11628 -2812
rect 11572 -2868 11574 -2822
rect 11574 -2868 11626 -2822
rect 11626 -2868 11628 -2822
rect 11572 -2938 11574 -2892
rect 11574 -2938 11626 -2892
rect 11626 -2938 11628 -2892
rect 11572 -2948 11628 -2938
rect 12832 -2822 12888 -2812
rect 12832 -2868 12834 -2822
rect 12834 -2868 12886 -2822
rect 12886 -2868 12888 -2822
rect 12832 -2938 12834 -2892
rect 12834 -2938 12886 -2892
rect 12886 -2938 12888 -2892
rect 12832 -2948 12888 -2938
rect 7864 -3159 7920 -3103
rect 10311 -3156 10313 -3134
rect 10313 -3156 10365 -3134
rect 10365 -3156 10367 -3134
rect 10311 -3168 10367 -3156
rect 10311 -3190 10313 -3168
rect 10313 -3190 10365 -3168
rect 10365 -3190 10367 -3168
rect 2052 -3938 2108 -3882
rect 2052 -4018 2108 -3962
rect 10311 -4159 10367 -4103
rect 7852 -4708 7908 -4652
rect 1912 -4824 1914 -4772
rect 1914 -4824 1966 -4772
rect 1966 -4824 1968 -4772
rect 1912 -4828 1968 -4824
rect 1912 -4888 1914 -4862
rect 1914 -4888 1966 -4862
rect 1966 -4888 1968 -4862
rect 1912 -4918 1968 -4888
rect 4912 -4848 4968 -4792
rect 6072 -4848 6128 -4792
rect 6152 -4848 6208 -4792
rect 6652 -4843 6708 -4787
rect 7472 -4843 7528 -4787
rect 8622 -4838 8678 -4782
rect 3762 -6111 3802 -6062
rect 3802 -6111 3818 -6062
rect 3852 -6111 3854 -6062
rect 3854 -6111 3866 -6062
rect 3866 -6111 3908 -6062
rect 3762 -6118 3818 -6111
rect 3852 -6118 3908 -6111
rect 5114 -6227 5170 -6225
rect 5194 -6227 5250 -6225
rect 5274 -6227 5330 -6225
rect 5354 -6227 5410 -6225
rect 5434 -6227 5490 -6225
rect 5514 -6227 5570 -6225
rect 5594 -6227 5650 -6225
rect 5674 -6227 5730 -6225
rect 5754 -6227 5810 -6225
rect 5834 -6227 5890 -6225
rect 5114 -6279 5124 -6227
rect 5124 -6279 5170 -6227
rect 5194 -6279 5240 -6227
rect 5240 -6279 5250 -6227
rect 5274 -6279 5304 -6227
rect 5304 -6279 5316 -6227
rect 5316 -6279 5330 -6227
rect 5354 -6279 5368 -6227
rect 5368 -6279 5380 -6227
rect 5380 -6279 5410 -6227
rect 5434 -6279 5444 -6227
rect 5444 -6279 5490 -6227
rect 5514 -6279 5560 -6227
rect 5560 -6279 5570 -6227
rect 5594 -6279 5624 -6227
rect 5624 -6279 5636 -6227
rect 5636 -6279 5650 -6227
rect 5674 -6279 5688 -6227
rect 5688 -6279 5700 -6227
rect 5700 -6279 5730 -6227
rect 5754 -6279 5764 -6227
rect 5764 -6279 5810 -6227
rect 5834 -6279 5880 -6227
rect 5880 -6279 5890 -6227
rect 5114 -6281 5170 -6279
rect 5194 -6281 5250 -6279
rect 5274 -6281 5330 -6279
rect 5354 -6281 5410 -6279
rect 5434 -6281 5490 -6279
rect 5514 -6281 5570 -6279
rect 5594 -6281 5650 -6279
rect 5674 -6281 5730 -6279
rect 5754 -6281 5810 -6279
rect 5834 -6281 5890 -6279
rect 4806 -6468 4862 -6458
rect 4806 -6514 4808 -6468
rect 4808 -6514 4860 -6468
rect 4860 -6514 4862 -6468
rect 4806 -6584 4808 -6538
rect 4808 -6584 4860 -6538
rect 4860 -6584 4862 -6538
rect 4806 -6594 4862 -6584
rect 6111 -6422 6113 -6376
rect 6113 -6422 6165 -6376
rect 6165 -6422 6167 -6376
rect 6111 -6432 6167 -6422
rect 6111 -6486 6113 -6456
rect 6113 -6486 6165 -6456
rect 6165 -6486 6167 -6456
rect 6111 -6498 6167 -6486
rect 6111 -6512 6113 -6498
rect 6113 -6512 6165 -6498
rect 6165 -6512 6167 -6498
rect 6111 -6550 6113 -6536
rect 6113 -6550 6165 -6536
rect 6165 -6550 6167 -6536
rect 6111 -6562 6167 -6550
rect 6111 -6592 6113 -6562
rect 6113 -6592 6165 -6562
rect 6165 -6592 6167 -6562
rect 6111 -6626 6167 -6616
rect 6111 -6672 6113 -6626
rect 6113 -6672 6165 -6626
rect 6165 -6672 6167 -6626
rect 7369 -6417 7371 -6371
rect 7371 -6417 7423 -6371
rect 7423 -6417 7425 -6371
rect 7369 -6427 7425 -6417
rect 7369 -6481 7371 -6451
rect 7371 -6481 7423 -6451
rect 7423 -6481 7425 -6451
rect 7369 -6493 7425 -6481
rect 7369 -6507 7371 -6493
rect 7371 -6507 7423 -6493
rect 7423 -6507 7425 -6493
rect 7369 -6545 7371 -6531
rect 7371 -6545 7423 -6531
rect 7423 -6545 7425 -6531
rect 7369 -6557 7425 -6545
rect 7369 -6587 7371 -6557
rect 7371 -6587 7423 -6557
rect 7423 -6587 7425 -6557
rect 7369 -6621 7425 -6611
rect 7369 -6667 7371 -6621
rect 7371 -6667 7423 -6621
rect 7423 -6667 7425 -6621
rect 6394 -6911 6450 -6909
rect 6474 -6911 6530 -6909
rect 6554 -6911 6610 -6909
rect 6634 -6911 6690 -6909
rect 6714 -6911 6770 -6909
rect 6794 -6911 6850 -6909
rect 6874 -6911 6930 -6909
rect 6954 -6911 7010 -6909
rect 7034 -6911 7090 -6909
rect 7114 -6911 7170 -6909
rect 6394 -6963 6404 -6911
rect 6404 -6963 6450 -6911
rect 6474 -6963 6520 -6911
rect 6520 -6963 6530 -6911
rect 6554 -6963 6584 -6911
rect 6584 -6963 6596 -6911
rect 6596 -6963 6610 -6911
rect 6634 -6963 6648 -6911
rect 6648 -6963 6660 -6911
rect 6660 -6963 6690 -6911
rect 6714 -6963 6724 -6911
rect 6724 -6963 6770 -6911
rect 6794 -6963 6840 -6911
rect 6840 -6963 6850 -6911
rect 6874 -6963 6904 -6911
rect 6904 -6963 6916 -6911
rect 6916 -6963 6930 -6911
rect 6954 -6963 6968 -6911
rect 6968 -6963 6980 -6911
rect 6980 -6963 7010 -6911
rect 7034 -6963 7044 -6911
rect 7044 -6963 7090 -6911
rect 7114 -6963 7160 -6911
rect 7160 -6963 7170 -6911
rect 6394 -6965 6450 -6963
rect 6474 -6965 6530 -6963
rect 6554 -6965 6610 -6963
rect 6634 -6965 6690 -6963
rect 6714 -6965 6770 -6963
rect 6794 -6965 6850 -6963
rect 6874 -6965 6930 -6963
rect 6954 -6965 7010 -6963
rect 7034 -6965 7090 -6963
rect 7114 -6965 7170 -6963
rect 8622 -7058 8678 -7032
rect 8622 -7088 8624 -7058
rect 8624 -7088 8676 -7058
rect 8676 -7088 8678 -7058
rect 8622 -7122 8678 -7112
rect 8622 -7168 8624 -7122
rect 8624 -7168 8676 -7122
rect 8676 -7168 8678 -7122
rect 8622 -7238 8624 -7192
rect 8624 -7238 8676 -7192
rect 8676 -7238 8678 -7192
rect 8622 -7248 8678 -7238
rect 8622 -7302 8624 -7272
rect 8624 -7302 8676 -7272
rect 8676 -7302 8678 -7272
rect 8622 -7328 8678 -7302
<< metal3 >>
rect 6540 128 6640 140
rect 6540 72 6562 128
rect 6618 72 6640 128
rect 6540 -682 6640 72
rect 10340 128 10420 140
rect 10340 72 10352 128
rect 10408 72 10420 128
rect 7630 -332 7730 -315
rect 7630 -388 7652 -332
rect 7708 -388 7730 -332
rect 7630 -412 7730 -388
rect 7630 -468 7652 -412
rect 7708 -468 7730 -412
rect 7630 -485 7730 -468
rect 2020 -748 2140 -720
rect 2020 -812 2048 -748
rect 2112 -812 2140 -748
rect 2020 -828 2140 -812
rect 2020 -892 2048 -828
rect 2112 -892 2140 -828
rect 2020 -1448 2140 -892
rect 3970 -748 4070 -735
rect 3970 -812 3988 -748
rect 4052 -812 4070 -748
rect 3970 -828 4070 -812
rect 3970 -892 3988 -828
rect 4052 -892 4070 -828
rect 3970 -905 4070 -892
rect 5230 -748 5330 -735
rect 5230 -812 5248 -748
rect 5312 -812 5330 -748
rect 5230 -828 5330 -812
rect 5230 -892 5248 -828
rect 5312 -892 5330 -828
rect 5230 -905 5330 -892
rect 6540 -738 6562 -682
rect 6618 -738 6640 -682
rect 10340 -700 10420 72
rect 6540 -762 6640 -738
rect 6540 -818 6562 -762
rect 6618 -818 6640 -762
rect 6540 -842 6640 -818
rect 6540 -898 6562 -842
rect 6618 -898 6640 -842
rect 6540 -922 6640 -898
rect 7750 -748 7850 -735
rect 7750 -812 7768 -748
rect 7832 -812 7850 -748
rect 7750 -828 7850 -812
rect 7750 -892 7768 -828
rect 7832 -892 7850 -828
rect 7750 -905 7850 -892
rect 9010 -748 9110 -735
rect 9010 -812 9028 -748
rect 9092 -812 9110 -748
rect 9010 -828 9110 -812
rect 9010 -892 9028 -828
rect 9092 -892 9110 -828
rect 9010 -905 9110 -892
rect 10340 -738 10422 -700
rect 10340 -794 10354 -738
rect 10410 -794 10422 -738
rect 10340 -818 10422 -794
rect 10340 -874 10354 -818
rect 10410 -874 10422 -818
rect 10340 -898 10422 -874
rect 6540 -978 6562 -922
rect 6618 -978 6640 -922
rect 6540 -1040 6640 -978
rect 10340 -954 10354 -898
rect 10410 -954 10422 -898
rect 11550 -748 11650 -735
rect 11550 -812 11568 -748
rect 11632 -812 11650 -748
rect 11550 -828 11650 -812
rect 11550 -892 11568 -828
rect 11632 -892 11650 -828
rect 11550 -905 11650 -892
rect 12810 -748 12910 -735
rect 12810 -812 12828 -748
rect 12892 -812 12910 -748
rect 12810 -828 12910 -812
rect 12810 -892 12828 -828
rect 12892 -892 12910 -828
rect 12810 -905 12910 -892
rect 10340 -991 10422 -954
rect 7820 -1059 7940 -1040
rect 7820 -1115 7853 -1059
rect 7909 -1115 7940 -1059
rect 2020 -1512 2048 -1448
rect 2112 -1512 2140 -1448
rect 2020 -1528 2140 -1512
rect 2020 -1592 2048 -1528
rect 2112 -1592 2140 -1528
rect 2020 -2148 2140 -1592
rect 3970 -1448 4070 -1435
rect 3970 -1512 3988 -1448
rect 4052 -1512 4070 -1448
rect 3970 -1528 4070 -1512
rect 3970 -1592 3988 -1528
rect 4052 -1592 4070 -1528
rect 3970 -1605 4070 -1592
rect 5250 -1448 5350 -1435
rect 5250 -1512 5268 -1448
rect 5332 -1512 5350 -1448
rect 5250 -1528 5350 -1512
rect 5250 -1592 5268 -1528
rect 5332 -1592 5350 -1528
rect 5250 -1605 5350 -1592
rect 6637 -1753 6728 -1720
rect 6637 -1809 6649 -1753
rect 6705 -1809 6728 -1753
rect 2020 -2212 2048 -2148
rect 2112 -2212 2140 -2148
rect 2020 -2228 2140 -2212
rect 2020 -2292 2048 -2228
rect 2112 -2292 2140 -2228
rect 2020 -2838 2140 -2292
rect 3970 -2148 4070 -2135
rect 3970 -2212 3988 -2148
rect 4052 -2212 4070 -2148
rect 3970 -2228 4070 -2212
rect 3970 -2292 3988 -2228
rect 4052 -2292 4070 -2228
rect 3970 -2305 4070 -2292
rect 5230 -2148 5330 -2135
rect 5230 -2212 5248 -2148
rect 5312 -2212 5330 -2148
rect 5230 -2228 5330 -2212
rect 5230 -2292 5248 -2228
rect 5312 -2292 5330 -2228
rect 5230 -2305 5330 -2292
rect 6637 -2434 6728 -1809
rect 6637 -2490 6651 -2434
rect 6707 -2490 6728 -2434
rect 2020 -2902 2048 -2838
rect 2112 -2902 2140 -2838
rect 2020 -3882 2140 -2902
rect 3970 -2808 4070 -2795
rect 3970 -2872 3988 -2808
rect 4052 -2872 4070 -2808
rect 3970 -2888 4070 -2872
rect 3970 -2952 3988 -2888
rect 4052 -2952 4070 -2888
rect 3970 -2965 4070 -2952
rect 5230 -2808 5330 -2795
rect 5230 -2872 5248 -2808
rect 5312 -2872 5330 -2808
rect 5230 -2888 5330 -2872
rect 5230 -2952 5248 -2888
rect 5312 -2952 5330 -2888
rect 5230 -2965 5330 -2952
rect 6637 -3080 6728 -2490
rect 6640 -3204 6728 -3080
rect 7820 -3094 7940 -1115
rect 10340 -1120 10420 -991
rect 9030 -1448 9130 -1435
rect 9030 -1512 9048 -1448
rect 9112 -1512 9130 -1448
rect 9030 -1528 9130 -1512
rect 9030 -1592 9048 -1528
rect 9112 -1592 9130 -1528
rect 9030 -1605 9130 -1592
rect 11550 -1448 11650 -1435
rect 11550 -1512 11568 -1448
rect 11632 -1512 11650 -1448
rect 11550 -1528 11650 -1512
rect 11550 -1592 11568 -1528
rect 11632 -1592 11650 -1528
rect 11550 -1605 11650 -1592
rect 12810 -1448 12910 -1435
rect 12810 -1512 12828 -1448
rect 12892 -1512 12910 -1448
rect 12810 -1528 12910 -1512
rect 12810 -1592 12828 -1528
rect 12892 -1592 12910 -1528
rect 12810 -1605 12910 -1592
rect 9030 -2148 9130 -2135
rect 9030 -2212 9048 -2148
rect 9112 -2212 9130 -2148
rect 9030 -2228 9130 -2212
rect 9030 -2292 9048 -2228
rect 9112 -2292 9130 -2228
rect 9030 -2305 9130 -2292
rect 11550 -2148 11650 -2135
rect 11550 -2212 11568 -2148
rect 11632 -2212 11650 -2148
rect 11550 -2228 11650 -2212
rect 11550 -2292 11568 -2228
rect 11632 -2292 11650 -2228
rect 11550 -2305 11650 -2292
rect 12810 -2148 12910 -2135
rect 12810 -2212 12828 -2148
rect 12892 -2212 12910 -2148
rect 12810 -2228 12910 -2212
rect 12810 -2292 12828 -2228
rect 12892 -2292 12910 -2228
rect 12810 -2305 12910 -2292
rect 9030 -2808 9130 -2795
rect 9030 -2872 9048 -2808
rect 9112 -2872 9130 -2808
rect 9030 -2888 9130 -2872
rect 9030 -2952 9048 -2888
rect 9112 -2952 9130 -2888
rect 9030 -2965 9130 -2952
rect 11550 -2808 11650 -2795
rect 11550 -2872 11568 -2808
rect 11632 -2872 11650 -2808
rect 11550 -2888 11650 -2872
rect 11550 -2952 11568 -2888
rect 11632 -2952 11650 -2888
rect 11550 -2965 11650 -2952
rect 12810 -2808 12910 -2795
rect 12810 -2872 12828 -2808
rect 12892 -2872 12910 -2808
rect 12810 -2888 12910 -2872
rect 12810 -2952 12828 -2888
rect 12892 -2952 12910 -2888
rect 12810 -2965 12910 -2952
rect 7820 -3103 7951 -3094
rect 7820 -3159 7864 -3103
rect 7920 -3159 7951 -3103
rect 7820 -3167 7951 -3159
rect 10298 -3134 10381 -3058
rect 6640 -3240 6724 -3204
rect 2020 -3938 2052 -3882
rect 2108 -3938 2140 -3882
rect 2020 -3962 2140 -3938
rect 2020 -4018 2052 -3962
rect 2108 -4018 2140 -3962
rect 2020 -4060 2140 -4018
rect 6636 -4640 6724 -3240
rect 1890 -4772 2010 -4740
rect 1890 -4828 1912 -4772
rect 1968 -4828 2010 -4772
rect 1890 -4862 2010 -4828
rect 1890 -4918 1912 -4862
rect 1968 -4918 2010 -4862
rect 1890 -6208 2010 -4918
rect 4890 -4792 4990 -4760
rect 4890 -4848 4912 -4792
rect 4968 -4848 4990 -4792
rect 4890 -5570 4990 -4848
rect 6030 -4792 6250 -4760
rect 6030 -4848 6072 -4792
rect 6128 -4848 6152 -4792
rect 6208 -4848 6250 -4792
rect 6030 -4880 6250 -4848
rect 6640 -4787 6720 -4640
rect 7820 -4652 7940 -3167
rect 10298 -3190 10311 -3134
rect 10367 -3190 10381 -3134
rect 10298 -4090 10381 -3190
rect 10298 -4103 10380 -4090
rect 10298 -4159 10311 -4103
rect 10367 -4159 10380 -4103
rect 10298 -4169 10380 -4159
rect 7820 -4708 7852 -4652
rect 7908 -4708 7940 -4652
rect 7820 -4720 7940 -4708
rect 6640 -4843 6652 -4787
rect 6708 -4843 6720 -4787
rect 6640 -4870 6720 -4843
rect 7460 -4787 7540 -4760
rect 7460 -4843 7472 -4787
rect 7528 -4843 7540 -4787
rect 7460 -4870 7540 -4843
rect 6090 -5570 6230 -4880
rect 7370 -4950 7540 -4870
rect 8590 -4782 8710 -4760
rect 8590 -4838 8622 -4782
rect 8678 -4838 8710 -4782
rect 7370 -5570 7450 -4950
rect 4888 -5630 4990 -5570
rect 6083 -5610 6230 -5570
rect 3750 -6048 3970 -6030
rect 3750 -6062 3768 -6048
rect 3832 -6062 3888 -6048
rect 3750 -6118 3762 -6062
rect 3832 -6112 3852 -6062
rect 3952 -6112 3970 -6048
rect 3818 -6118 3852 -6112
rect 3908 -6118 3970 -6112
rect 3750 -6130 3970 -6118
rect 1890 -6272 1918 -6208
rect 1982 -6272 2010 -6208
rect 1890 -6848 2010 -6272
rect 4888 -6308 4985 -5630
rect 5100 -6221 5905 -6215
rect 5100 -6285 5110 -6221
rect 5174 -6285 5190 -6221
rect 5254 -6285 5270 -6221
rect 5334 -6285 5350 -6221
rect 5414 -6285 5430 -6221
rect 5494 -6285 5510 -6221
rect 5574 -6285 5590 -6221
rect 5654 -6285 5670 -6221
rect 5734 -6285 5750 -6221
rect 5814 -6285 5830 -6221
rect 5894 -6285 5905 -6221
rect 5100 -6291 5905 -6285
rect 4796 -6433 4985 -6308
rect 4790 -6458 4985 -6433
rect 4790 -6514 4806 -6458
rect 4862 -6514 4985 -6458
rect 4790 -6538 4985 -6514
rect 4790 -6594 4806 -6538
rect 4862 -6594 4985 -6538
rect 4790 -6618 4985 -6594
rect 4791 -6702 4985 -6618
rect 4846 -6711 4985 -6702
rect 6083 -6376 6227 -5610
rect 7357 -6357 7454 -5570
rect 6083 -6432 6111 -6376
rect 6167 -6432 6227 -6376
rect 6083 -6456 6227 -6432
rect 6083 -6512 6111 -6456
rect 6167 -6512 6227 -6456
rect 6083 -6536 6227 -6512
rect 6083 -6592 6111 -6536
rect 6167 -6592 6227 -6536
rect 6083 -6616 6227 -6592
rect 6083 -6672 6111 -6616
rect 6167 -6672 6227 -6616
rect 4846 -6722 4955 -6711
rect 6083 -6716 6227 -6672
rect 7352 -6371 7454 -6357
rect 7352 -6427 7369 -6371
rect 7425 -6427 7454 -6371
rect 7352 -6451 7454 -6427
rect 7352 -6507 7369 -6451
rect 7425 -6507 7454 -6451
rect 7352 -6531 7454 -6507
rect 7352 -6587 7369 -6531
rect 7425 -6587 7454 -6531
rect 7352 -6611 7454 -6587
rect 7352 -6667 7369 -6611
rect 7425 -6667 7454 -6611
rect 7352 -6680 7454 -6667
rect 7357 -6697 7454 -6680
rect 1890 -6912 1918 -6848
rect 1982 -6912 2010 -6848
rect 1890 -6930 2010 -6912
rect 6380 -6905 7185 -6899
rect 6380 -6969 6390 -6905
rect 6454 -6969 6470 -6905
rect 6534 -6969 6550 -6905
rect 6614 -6969 6630 -6905
rect 6694 -6969 6710 -6905
rect 6774 -6969 6790 -6905
rect 6854 -6969 6870 -6905
rect 6934 -6969 6950 -6905
rect 7014 -6969 7030 -6905
rect 7094 -6969 7110 -6905
rect 7174 -6969 7185 -6905
rect 6380 -6975 7185 -6969
rect 8590 -7032 8710 -4838
rect 8590 -7088 8622 -7032
rect 8678 -7088 8710 -7032
rect 8590 -7112 8710 -7088
rect 8590 -7168 8622 -7112
rect 8678 -7168 8710 -7112
rect 8590 -7192 8710 -7168
rect 8590 -7248 8622 -7192
rect 8678 -7248 8710 -7192
rect 8590 -7272 8710 -7248
rect 8590 -7328 8622 -7272
rect 8678 -7328 8710 -7272
rect 8590 -7390 8710 -7328
<< via3 >>
rect 2048 -812 2112 -748
rect 2048 -892 2112 -828
rect 3988 -752 4052 -748
rect 3988 -808 3992 -752
rect 3992 -808 4048 -752
rect 4048 -808 4052 -752
rect 3988 -812 4052 -808
rect 3988 -832 4052 -828
rect 3988 -888 3992 -832
rect 3992 -888 4048 -832
rect 4048 -888 4052 -832
rect 3988 -892 4052 -888
rect 5248 -752 5312 -748
rect 5248 -808 5252 -752
rect 5252 -808 5308 -752
rect 5308 -808 5312 -752
rect 5248 -812 5312 -808
rect 5248 -832 5312 -828
rect 5248 -888 5252 -832
rect 5252 -888 5308 -832
rect 5308 -888 5312 -832
rect 5248 -892 5312 -888
rect 7768 -752 7832 -748
rect 7768 -808 7772 -752
rect 7772 -808 7828 -752
rect 7828 -808 7832 -752
rect 7768 -812 7832 -808
rect 7768 -832 7832 -828
rect 7768 -888 7772 -832
rect 7772 -888 7828 -832
rect 7828 -888 7832 -832
rect 7768 -892 7832 -888
rect 9028 -752 9092 -748
rect 9028 -808 9032 -752
rect 9032 -808 9088 -752
rect 9088 -808 9092 -752
rect 9028 -812 9092 -808
rect 9028 -832 9092 -828
rect 9028 -888 9032 -832
rect 9032 -888 9088 -832
rect 9088 -888 9092 -832
rect 9028 -892 9092 -888
rect 11568 -752 11632 -748
rect 11568 -808 11572 -752
rect 11572 -808 11628 -752
rect 11628 -808 11632 -752
rect 11568 -812 11632 -808
rect 11568 -832 11632 -828
rect 11568 -888 11572 -832
rect 11572 -888 11628 -832
rect 11628 -888 11632 -832
rect 11568 -892 11632 -888
rect 12828 -752 12892 -748
rect 12828 -808 12832 -752
rect 12832 -808 12888 -752
rect 12888 -808 12892 -752
rect 12828 -812 12892 -808
rect 12828 -832 12892 -828
rect 12828 -888 12832 -832
rect 12832 -888 12888 -832
rect 12888 -888 12892 -832
rect 12828 -892 12892 -888
rect 2048 -1512 2112 -1448
rect 2048 -1592 2112 -1528
rect 3988 -1452 4052 -1448
rect 3988 -1508 3992 -1452
rect 3992 -1508 4048 -1452
rect 4048 -1508 4052 -1452
rect 3988 -1512 4052 -1508
rect 3988 -1532 4052 -1528
rect 3988 -1588 3992 -1532
rect 3992 -1588 4048 -1532
rect 4048 -1588 4052 -1532
rect 3988 -1592 4052 -1588
rect 5268 -1452 5332 -1448
rect 5268 -1508 5272 -1452
rect 5272 -1508 5328 -1452
rect 5328 -1508 5332 -1452
rect 5268 -1512 5332 -1508
rect 5268 -1532 5332 -1528
rect 5268 -1588 5272 -1532
rect 5272 -1588 5328 -1532
rect 5328 -1588 5332 -1532
rect 5268 -1592 5332 -1588
rect 2048 -2212 2112 -2148
rect 2048 -2292 2112 -2228
rect 3988 -2152 4052 -2148
rect 3988 -2208 3992 -2152
rect 3992 -2208 4048 -2152
rect 4048 -2208 4052 -2152
rect 3988 -2212 4052 -2208
rect 3988 -2232 4052 -2228
rect 3988 -2288 3992 -2232
rect 3992 -2288 4048 -2232
rect 4048 -2288 4052 -2232
rect 3988 -2292 4052 -2288
rect 5248 -2152 5312 -2148
rect 5248 -2208 5252 -2152
rect 5252 -2208 5308 -2152
rect 5308 -2208 5312 -2152
rect 5248 -2212 5312 -2208
rect 5248 -2232 5312 -2228
rect 5248 -2288 5252 -2232
rect 5252 -2288 5308 -2232
rect 5308 -2288 5312 -2232
rect 5248 -2292 5312 -2288
rect 2048 -2902 2112 -2838
rect 3988 -2812 4052 -2808
rect 3988 -2868 3992 -2812
rect 3992 -2868 4048 -2812
rect 4048 -2868 4052 -2812
rect 3988 -2872 4052 -2868
rect 3988 -2892 4052 -2888
rect 3988 -2948 3992 -2892
rect 3992 -2948 4048 -2892
rect 4048 -2948 4052 -2892
rect 3988 -2952 4052 -2948
rect 5248 -2812 5312 -2808
rect 5248 -2868 5252 -2812
rect 5252 -2868 5308 -2812
rect 5308 -2868 5312 -2812
rect 5248 -2872 5312 -2868
rect 5248 -2892 5312 -2888
rect 5248 -2948 5252 -2892
rect 5252 -2948 5308 -2892
rect 5308 -2948 5312 -2892
rect 5248 -2952 5312 -2948
rect 9048 -1452 9112 -1448
rect 9048 -1508 9052 -1452
rect 9052 -1508 9108 -1452
rect 9108 -1508 9112 -1452
rect 9048 -1512 9112 -1508
rect 9048 -1532 9112 -1528
rect 9048 -1588 9052 -1532
rect 9052 -1588 9108 -1532
rect 9108 -1588 9112 -1532
rect 9048 -1592 9112 -1588
rect 11568 -1452 11632 -1448
rect 11568 -1508 11572 -1452
rect 11572 -1508 11628 -1452
rect 11628 -1508 11632 -1452
rect 11568 -1512 11632 -1508
rect 11568 -1532 11632 -1528
rect 11568 -1588 11572 -1532
rect 11572 -1588 11628 -1532
rect 11628 -1588 11632 -1532
rect 11568 -1592 11632 -1588
rect 12828 -1452 12892 -1448
rect 12828 -1508 12832 -1452
rect 12832 -1508 12888 -1452
rect 12888 -1508 12892 -1452
rect 12828 -1512 12892 -1508
rect 12828 -1532 12892 -1528
rect 12828 -1588 12832 -1532
rect 12832 -1588 12888 -1532
rect 12888 -1588 12892 -1532
rect 12828 -1592 12892 -1588
rect 9048 -2152 9112 -2148
rect 9048 -2208 9052 -2152
rect 9052 -2208 9108 -2152
rect 9108 -2208 9112 -2152
rect 9048 -2212 9112 -2208
rect 9048 -2232 9112 -2228
rect 9048 -2288 9052 -2232
rect 9052 -2288 9108 -2232
rect 9108 -2288 9112 -2232
rect 9048 -2292 9112 -2288
rect 11568 -2152 11632 -2148
rect 11568 -2208 11572 -2152
rect 11572 -2208 11628 -2152
rect 11628 -2208 11632 -2152
rect 11568 -2212 11632 -2208
rect 11568 -2232 11632 -2228
rect 11568 -2288 11572 -2232
rect 11572 -2288 11628 -2232
rect 11628 -2288 11632 -2232
rect 11568 -2292 11632 -2288
rect 12828 -2152 12892 -2148
rect 12828 -2208 12832 -2152
rect 12832 -2208 12888 -2152
rect 12888 -2208 12892 -2152
rect 12828 -2212 12892 -2208
rect 12828 -2232 12892 -2228
rect 12828 -2288 12832 -2232
rect 12832 -2288 12888 -2232
rect 12888 -2288 12892 -2232
rect 12828 -2292 12892 -2288
rect 9048 -2812 9112 -2808
rect 9048 -2868 9052 -2812
rect 9052 -2868 9108 -2812
rect 9108 -2868 9112 -2812
rect 9048 -2872 9112 -2868
rect 9048 -2892 9112 -2888
rect 9048 -2948 9052 -2892
rect 9052 -2948 9108 -2892
rect 9108 -2948 9112 -2892
rect 9048 -2952 9112 -2948
rect 11568 -2812 11632 -2808
rect 11568 -2868 11572 -2812
rect 11572 -2868 11628 -2812
rect 11628 -2868 11632 -2812
rect 11568 -2872 11632 -2868
rect 11568 -2892 11632 -2888
rect 11568 -2948 11572 -2892
rect 11572 -2948 11628 -2892
rect 11628 -2948 11632 -2892
rect 11568 -2952 11632 -2948
rect 12828 -2812 12892 -2808
rect 12828 -2868 12832 -2812
rect 12832 -2868 12888 -2812
rect 12888 -2868 12892 -2812
rect 12828 -2872 12892 -2868
rect 12828 -2892 12892 -2888
rect 12828 -2948 12832 -2892
rect 12832 -2948 12888 -2892
rect 12888 -2948 12892 -2892
rect 12828 -2952 12892 -2948
rect 3768 -6062 3832 -6048
rect 3888 -6062 3952 -6048
rect 3768 -6112 3818 -6062
rect 3818 -6112 3832 -6062
rect 3888 -6112 3908 -6062
rect 3908 -6112 3952 -6062
rect 1918 -6272 1982 -6208
rect 5110 -6225 5174 -6221
rect 5110 -6281 5114 -6225
rect 5114 -6281 5170 -6225
rect 5170 -6281 5174 -6225
rect 5110 -6285 5174 -6281
rect 5190 -6225 5254 -6221
rect 5190 -6281 5194 -6225
rect 5194 -6281 5250 -6225
rect 5250 -6281 5254 -6225
rect 5190 -6285 5254 -6281
rect 5270 -6225 5334 -6221
rect 5270 -6281 5274 -6225
rect 5274 -6281 5330 -6225
rect 5330 -6281 5334 -6225
rect 5270 -6285 5334 -6281
rect 5350 -6225 5414 -6221
rect 5350 -6281 5354 -6225
rect 5354 -6281 5410 -6225
rect 5410 -6281 5414 -6225
rect 5350 -6285 5414 -6281
rect 5430 -6225 5494 -6221
rect 5430 -6281 5434 -6225
rect 5434 -6281 5490 -6225
rect 5490 -6281 5494 -6225
rect 5430 -6285 5494 -6281
rect 5510 -6225 5574 -6221
rect 5510 -6281 5514 -6225
rect 5514 -6281 5570 -6225
rect 5570 -6281 5574 -6225
rect 5510 -6285 5574 -6281
rect 5590 -6225 5654 -6221
rect 5590 -6281 5594 -6225
rect 5594 -6281 5650 -6225
rect 5650 -6281 5654 -6225
rect 5590 -6285 5654 -6281
rect 5670 -6225 5734 -6221
rect 5670 -6281 5674 -6225
rect 5674 -6281 5730 -6225
rect 5730 -6281 5734 -6225
rect 5670 -6285 5734 -6281
rect 5750 -6225 5814 -6221
rect 5750 -6281 5754 -6225
rect 5754 -6281 5810 -6225
rect 5810 -6281 5814 -6225
rect 5750 -6285 5814 -6281
rect 5830 -6225 5894 -6221
rect 5830 -6281 5834 -6225
rect 5834 -6281 5890 -6225
rect 5890 -6281 5894 -6225
rect 5830 -6285 5894 -6281
rect 1918 -6912 1982 -6848
rect 6390 -6909 6454 -6905
rect 6390 -6965 6394 -6909
rect 6394 -6965 6450 -6909
rect 6450 -6965 6454 -6909
rect 6390 -6969 6454 -6965
rect 6470 -6909 6534 -6905
rect 6470 -6965 6474 -6909
rect 6474 -6965 6530 -6909
rect 6530 -6965 6534 -6909
rect 6470 -6969 6534 -6965
rect 6550 -6909 6614 -6905
rect 6550 -6965 6554 -6909
rect 6554 -6965 6610 -6909
rect 6610 -6965 6614 -6909
rect 6550 -6969 6614 -6965
rect 6630 -6909 6694 -6905
rect 6630 -6965 6634 -6909
rect 6634 -6965 6690 -6909
rect 6690 -6965 6694 -6909
rect 6630 -6969 6694 -6965
rect 6710 -6909 6774 -6905
rect 6710 -6965 6714 -6909
rect 6714 -6965 6770 -6909
rect 6770 -6965 6774 -6909
rect 6710 -6969 6774 -6965
rect 6790 -6909 6854 -6905
rect 6790 -6965 6794 -6909
rect 6794 -6965 6850 -6909
rect 6850 -6965 6854 -6909
rect 6790 -6969 6854 -6965
rect 6870 -6909 6934 -6905
rect 6870 -6965 6874 -6909
rect 6874 -6965 6930 -6909
rect 6930 -6965 6934 -6909
rect 6870 -6969 6934 -6965
rect 6950 -6909 7014 -6905
rect 6950 -6965 6954 -6909
rect 6954 -6965 7010 -6909
rect 7010 -6965 7014 -6909
rect 6950 -6969 7014 -6965
rect 7030 -6909 7094 -6905
rect 7030 -6965 7034 -6909
rect 7034 -6965 7090 -6909
rect 7090 -6965 7094 -6909
rect 7030 -6969 7094 -6965
rect 7110 -6909 7174 -6905
rect 7110 -6965 7114 -6909
rect 7114 -6965 7170 -6909
rect 7170 -6965 7174 -6909
rect 7110 -6969 7174 -6965
<< metal4 >>
rect 2020 -739 12900 -720
rect 2020 -748 12901 -739
rect 2020 -812 2048 -748
rect 2112 -812 3988 -748
rect 4052 -812 5248 -748
rect 5312 -812 7768 -748
rect 7832 -812 9028 -748
rect 9092 -812 11568 -748
rect 11632 -812 12828 -748
rect 12892 -812 12901 -748
rect 2020 -828 12901 -812
rect 2020 -892 2048 -828
rect 2112 -892 3988 -828
rect 4052 -892 5248 -828
rect 5312 -892 7768 -828
rect 7832 -892 9028 -828
rect 9092 -892 11568 -828
rect 11632 -892 12828 -828
rect 12892 -892 12901 -828
rect 2020 -901 12901 -892
rect 2020 -920 12900 -901
rect 2020 -1439 12900 -1420
rect 2020 -1448 12901 -1439
rect 2020 -1512 2048 -1448
rect 2112 -1512 3988 -1448
rect 4052 -1512 5268 -1448
rect 5332 -1512 9048 -1448
rect 9112 -1512 11568 -1448
rect 11632 -1512 12828 -1448
rect 12892 -1512 12901 -1448
rect 2020 -1528 12901 -1512
rect 2020 -1592 2048 -1528
rect 2112 -1592 3988 -1528
rect 4052 -1592 5268 -1528
rect 5332 -1592 9048 -1528
rect 9112 -1592 11568 -1528
rect 11632 -1592 12828 -1528
rect 12892 -1592 12901 -1528
rect 2020 -1600 12901 -1592
rect 2020 -1620 7720 -1600
rect 8200 -1601 12901 -1600
rect 8200 -1620 12900 -1601
rect 2020 -2139 12900 -2120
rect 2020 -2148 12901 -2139
rect 2020 -2212 2048 -2148
rect 2112 -2212 3988 -2148
rect 4052 -2212 5248 -2148
rect 5312 -2212 9048 -2148
rect 9112 -2212 11568 -2148
rect 11632 -2212 12828 -2148
rect 12892 -2212 12901 -2148
rect 2020 -2228 12901 -2212
rect 2020 -2292 2048 -2228
rect 2112 -2292 3988 -2228
rect 4052 -2292 5248 -2228
rect 5312 -2292 9048 -2228
rect 9112 -2292 11568 -2228
rect 11632 -2292 12828 -2228
rect 12892 -2292 12901 -2228
rect 2020 -2301 12901 -2292
rect 2020 -2320 12900 -2301
rect 2020 -2780 7740 -2771
rect 8060 -2780 12904 -2771
rect 2020 -2808 12904 -2780
rect 2020 -2838 3988 -2808
rect 2020 -2902 2048 -2838
rect 2112 -2872 3988 -2838
rect 4052 -2872 5248 -2808
rect 5312 -2872 9048 -2808
rect 9112 -2872 11568 -2808
rect 11632 -2872 12828 -2808
rect 12892 -2872 12904 -2808
rect 2112 -2888 12904 -2872
rect 2112 -2902 3988 -2888
rect 2020 -2952 3988 -2902
rect 4052 -2952 5248 -2888
rect 5312 -2952 9048 -2888
rect 9112 -2952 11568 -2888
rect 11632 -2952 12828 -2888
rect 12892 -2952 12904 -2888
rect 2020 -2960 12904 -2952
rect 2020 -2971 7740 -2960
rect 8060 -2971 12904 -2960
rect 2020 -4070 2140 -3790
rect 3750 -6048 3970 -6030
rect 3750 -6050 3768 -6048
rect 1820 -6112 3768 -6050
rect 3832 -6112 3888 -6048
rect 3952 -6112 3970 -6048
rect 1820 -6130 3970 -6112
rect 1890 -6208 6010 -6190
rect 1890 -6272 1918 -6208
rect 1982 -6221 6010 -6208
rect 1982 -6270 5110 -6221
rect 1982 -6272 2010 -6270
rect 1890 -6290 2010 -6272
rect 4990 -6285 5110 -6270
rect 5174 -6285 5190 -6221
rect 5254 -6285 5270 -6221
rect 5334 -6285 5350 -6221
rect 5414 -6285 5430 -6221
rect 5494 -6285 5510 -6221
rect 5574 -6285 5590 -6221
rect 5654 -6285 5670 -6221
rect 5734 -6285 5750 -6221
rect 5814 -6285 5830 -6221
rect 5894 -6285 6010 -6221
rect 4990 -6310 6010 -6285
rect 1890 -6848 2010 -6830
rect 1890 -6912 1918 -6848
rect 1982 -6870 2010 -6848
rect 3060 -6870 3750 -6850
rect 1982 -6905 7250 -6870
rect 1982 -6912 6390 -6905
rect 1890 -6930 6390 -6912
rect 6230 -6969 6390 -6930
rect 6454 -6969 6470 -6905
rect 6534 -6969 6550 -6905
rect 6614 -6969 6630 -6905
rect 6694 -6969 6710 -6905
rect 6774 -6969 6790 -6905
rect 6854 -6969 6870 -6905
rect 6934 -6969 6950 -6905
rect 7014 -6969 7030 -6905
rect 7094 -6969 7110 -6905
rect 7174 -6969 7250 -6905
rect 6230 -6990 7250 -6969
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M32_A
timestamp 1757161594
transform 0 1 7250 -1 0 -1510
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M32_B
timestamp 1757161594
transform 0 1 8512 -1 0 -1510
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M32_C
timestamp 1757161594
transform 0 1 7250 -1 0 -2196
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M32_D
timestamp 1757161594
transform 0 1 8512 -1 0 -2196
box -396 -684 396 684
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M33_A
timestamp 1757161594
transform 0 1 5530 -1 0 -7193
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M33_B
timestamp 1757161594
transform 0 1 6790 -1 0 -6513
box -386 -669 386 669
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M34_A
timestamp 1757161594
transform 0 1 7250 -1 0 -824
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M34_B
timestamp 1757161594
transform 0 1 8512 -1 0 -824
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M34_C
timestamp 1757161594
transform 0 1 7250 -1 0 -2882
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M34_D
timestamp 1757161594
transform 0 1 8512 -1 0 -2882
box -396 -684 396 684
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M35_A
timestamp 1757161594
transform 0 1 4289 -1 0 -5834
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M35_B
timestamp 1757161594
transform 0 1 5540 -1 0 -5834
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M35_C
timestamp 1757161594
transform 0 1 6789 -1 0 -5834
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M35_D
timestamp 1757161594
transform 0 1 8030 -1 0 -5833
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M35_E
timestamp 1757161594
transform 0 1 4290 -1 0 -7873
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M35_F
timestamp 1757161594
transform 0 1 5530 -1 0 -7873
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M35_G
timestamp 1757161594
transform 0 1 6770 -1 0 -7873
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M36_A
timestamp 1757161594
transform 0 1 4289 -1 0 -7194
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M36_B
timestamp 1757161594
transform 0 1 8029 -1 0 -6514
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M37_A
timestamp 1757161594
transform 0 1 4290 -1 0 -6513
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M37_B
timestamp 1757161594
transform 0 1 8030 -1 0 -7193
box -386 -669 386 669
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M38_A
timestamp 1757161594
transform 0 1 5988 -1 0 -824
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M38_B
timestamp 1757161594
transform 0 1 5988 -1 0 -2882
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M38_C
timestamp 1757161594
transform 0 1 9774 -1 0 -824
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M38_D
timestamp 1757161594
transform 0 1 9774 -1 0 -2882
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M39_A
timestamp 1757161594
transform 0 1 5988 -1 0 -1510
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M39_B
timestamp 1757161594
transform 0 1 5988 -1 0 -2196
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M39_C
timestamp 1757161594
transform 0 1 9774 -1 0 -1510
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M39_D
timestamp 1757161594
transform 0 1 9774 -1 0 -2196
box -396 -684 396 684
use sky130_fd_pr__nfet_01v8_lvt_PAU7SL  M40
timestamp 1757161594
transform 0 1 2269 -1 0 -4844
box -286 -369 286 369
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M41_A
timestamp 1757161594
transform 0 1 5530 -1 0 -6513
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  M41_B
timestamp 1757161594
transform 0 1 6770 -1 0 -7193
box -386 -669 386 669
use sky130_fd_pr__pfet_01v8_lvt_9UXMRD  M42_A
timestamp 1757161594
transform 1 0 4196 0 1 464
box -2196 -284 2196 284
use sky130_fd_pr__pfet_01v8_lvt_LVXMRT  M42_B
timestamp 1757161594
transform 1 0 8482 0 1 464
box -2196 -284 2196 284
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M43_1
timestamp 1757161594
transform 0 1 3464 -1 0 -824
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M43_2
timestamp 1757161594
transform 0 1 4726 -1 0 -824
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M43_3
timestamp 1757161594
transform 0 1 11036 -1 0 -2882
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M43_4
timestamp 1757161594
transform 0 1 12298 -1 0 -2882
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M44_1
timestamp 1757161594
transform 0 1 3464 -1 0 -1510
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M44_2
timestamp 1757161594
transform 0 1 4726 -1 0 -1510
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M44_3
timestamp 1757161594
transform 0 1 11036 -1 0 -2196
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M44_4
timestamp 1757161594
transform 0 1 12298 -1 0 -2196
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M45_1
timestamp 1757161594
transform 0 1 3464 -1 0 -2196
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M45_2
timestamp 1757161594
transform 0 1 4726 -1 0 -2196
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M45_3
timestamp 1757161594
transform 0 1 11036 -1 0 -1510
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M45_4
timestamp 1757161594
transform 0 1 12298 -1 0 -1510
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M46_2
timestamp 1757161594
transform 0 1 7244 -1 0 -3564
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M46_3
timestamp 1757161594
transform 0 1 11036 -1 0 -824
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  M46_4
timestamp 1757161594
transform 0 1 12298 -1 0 -824
box -396 -684 396 684
use sky130_fd_pr__nfet_01v8_lvt_V2BN2G  sky130_fd_pr__nfet_01v8_lvt_V2BN2G_0
timestamp 1757161594
transform 0 1 3340 -1 0 -8563
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_0
timestamp 1757161594
transform 0 1 3339 -1 0 -7194
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_1
timestamp 1757161594
transform 0 1 8981 -1 0 -7191
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_2
timestamp 1757161594
transform 0 1 3339 -1 0 -7875
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_3
timestamp 1757161594
transform 0 1 3339 -1 0 -6508
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_4
timestamp 1757161594
transform 0 1 3338 -1 0 -5834
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_5
timestamp 1757161594
transform 0 1 3338 -1 0 -5149
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_7
timestamp 1757161594
transform 0 1 8982 -1 0 -8564
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_8
timestamp 1757161594
transform 0 1 8981 -1 0 -7873
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_9
timestamp 1757161594
transform 0 1 8982 -1 0 -6514
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_10
timestamp 1757161594
transform 0 1 8983 -1 0 -5833
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_VYCASF  sky130_fd_pr__nfet_01v8_lvt_VYCASF_11
timestamp 1757161594
transform 0 1 8983 -1 0 -5151
box -386 -369 386 369
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_0
timestamp 1757161594
transform 0 1 8030 -1 0 -7873
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_1
timestamp 1757161594
transform 0 1 8029 -1 0 -8564
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_2
timestamp 1757161594
transform 0 1 4291 -1 0 -8562
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_3
timestamp 1757161594
transform 0 1 5534 -1 0 -8562
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_4
timestamp 1757161594
transform 0 1 6773 -1 0 -8563
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_5
timestamp 1757161594
transform 0 1 6794 -1 0 -5148
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_6
timestamp 1757161594
transform 0 1 5541 -1 0 -5148
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_7
timestamp 1757161594
transform 0 1 4290 -1 0 -5150
box -386 -669 386 669
use sky130_fd_pr__nfet_01v8_lvt_ZVWESF  sky130_fd_pr__nfet_01v8_lvt_ZVWESF_8
timestamp 1757161594
transform 0 1 8028 -1 0 -5149
box -386 -669 386 669
use sky130_fd_pr__pfet_01v8_lvt_2QSR6E  sky130_fd_pr__pfet_01v8_lvt_2QSR6E_0
timestamp 1757161594
transform 0 1 13264 -1 0 -144
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_0
timestamp 1757161594
transform 0 1 2504 -1 0 -3564
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_1
timestamp 1757161594
transform 0 1 13264 -1 0 -2884
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_2
timestamp 1757161594
transform 0 1 13264 -1 0 -2204
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_3
timestamp 1757161594
transform 0 1 13264 -1 0 -1524
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_5
timestamp 1757161594
transform 0 1 13264 -1 0 -844
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_6
timestamp 1757161594
transform 0 1 13264 -1 0 -3564
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_7
timestamp 1757161594
transform 0 1 2504 -1 0 -2884
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_8
timestamp 1757161594
transform 0 1 2504 -1 0 -2204
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_9
timestamp 1757161594
transform 0 1 2504 -1 0 -1524
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_10
timestamp 1757161594
transform 0 1 2504 -1 0 -144
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_JY4D7E  sky130_fd_pr__pfet_01v8_lvt_JY4D7E_11
timestamp 1757161594
transform 0 1 2504 -1 0 -824
box -396 -384 396 384
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_0
timestamp 1757161594
transform 0 1 3464 -1 0 -2882
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_1
timestamp 1757161594
transform 0 1 4726 -1 0 -2882
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_3
timestamp 1757161594
transform 0 1 4724 -1 0 -3564
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_4
timestamp 1757161594
transform 0 1 5984 -1 0 -3564
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_5
timestamp 1757161594
transform 0 1 11029 -1 0 -3564
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_6
timestamp 1757161594
transform 0 1 8504 -1 0 -3564
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_7
timestamp 1757161594
transform 0 1 9764 -1 0 -3564
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_8
timestamp 1757161594
transform 0 1 12298 -1 0 -3564
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_9
timestamp 1757161594
transform 0 1 12299 -1 0 -144
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_10
timestamp 1757161594
transform 0 1 3464 -1 0 -144
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_11
timestamp 1757161594
transform 0 1 4724 -1 0 -144
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_12
timestamp 1757161594
transform 0 1 5984 -1 0 -144
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_13
timestamp 1757161594
transform 0 1 7244 -1 0 -144
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_14
timestamp 1757161594
transform 0 1 8504 -1 0 -144
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_15
timestamp 1757161594
transform 0 1 9764 -1 0 -144
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_NVX44G  sky130_fd_pr__pfet_01v8_lvt_NVX44G_16
timestamp 1757161594
transform 0 1 11024 -1 0 -144
box -396 -684 396 684
use sky130_fd_pr__pfet_01v8_lvt_UY454G  sky130_fd_pr__pfet_01v8_lvt_UY454G_0
timestamp 1757161594
transform 0 1 3464 -1 0 -3564
box -396 -684 396 684
<< labels >>
rlabel metal2 s 3940 -3960 4020 -3880 4 PBias
port 0 nsew
rlabel metal2 s 13880 -4280 13960 -4200 4 Vbias1
port 1 nsew
rlabel metal2 s 13880 -4390 13960 -4310 4 Vbias2
port 2 nsew
rlabel metal2 s 13880 -4500 13960 -4420 4 Vbias3
port 3 nsew
rlabel metal2 s 13880 -4610 13960 -4530 4 Vbias4
port 4 nsew
<< end >>
