magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect 60 3020 280 3030
rect -290 2380 4270 3020
rect -290 2320 3680 2380
rect 3860 2320 4270 2380
rect -290 -530 4270 2320
<< nsubdiff >>
rect -247 2883 -185 2917
rect -151 2883 -117 2917
rect -83 2883 -49 2917
rect -15 2883 19 2917
rect 53 2883 87 2917
rect 121 2883 155 2917
rect 189 2883 223 2917
rect 257 2883 291 2917
rect 325 2883 359 2917
rect 393 2883 427 2917
rect 461 2883 495 2917
rect 529 2883 563 2917
rect 597 2883 631 2917
rect 665 2883 699 2917
rect 733 2883 767 2917
rect 801 2883 835 2917
rect 869 2883 903 2917
rect 937 2883 971 2917
rect 1005 2883 1039 2917
rect 1073 2883 1107 2917
rect 1141 2883 1175 2917
rect 1209 2883 1243 2917
rect 1277 2883 1311 2917
rect 1345 2883 1379 2917
rect 1413 2883 1447 2917
rect 1481 2883 1515 2917
rect 1549 2883 1583 2917
rect 1617 2883 1651 2917
rect 1685 2883 1719 2917
rect 1753 2883 1787 2917
rect 1821 2883 1855 2917
rect 1889 2883 1923 2917
rect 1957 2883 1991 2917
rect 2025 2883 2059 2917
rect 2093 2883 2127 2917
rect 2161 2883 2195 2917
rect 2229 2883 2263 2917
rect 2297 2883 2331 2917
rect 2365 2883 2399 2917
rect 2433 2883 2467 2917
rect 2501 2883 2535 2917
rect 2569 2883 2603 2917
rect 2637 2883 2671 2917
rect 2705 2883 2739 2917
rect 2773 2883 2807 2917
rect 2841 2883 2875 2917
rect 2909 2883 2943 2917
rect 2977 2883 3011 2917
rect 3045 2883 3079 2917
rect 3113 2883 3147 2917
rect 3181 2883 3215 2917
rect 3249 2883 3283 2917
rect 3317 2883 3351 2917
rect 3385 2883 3419 2917
rect 3453 2883 3487 2917
rect 3521 2883 3555 2917
rect 3589 2883 3623 2917
rect 3657 2883 3691 2917
rect 3725 2883 3759 2917
rect 3793 2883 3827 2917
rect 3861 2883 3895 2917
rect 3929 2883 3963 2917
rect 3997 2883 4031 2917
rect 4065 2883 4127 2917
rect -247 2835 -213 2883
rect -247 2767 -213 2801
rect -247 2699 -213 2733
rect -247 2631 -213 2665
rect -247 2563 -213 2597
rect -247 2495 -213 2529
rect -247 2427 -213 2461
rect -247 2359 -213 2393
rect -247 2291 -213 2325
rect -247 2223 -213 2257
rect -247 2155 -213 2189
rect -247 2087 -213 2121
rect -247 2019 -213 2053
rect -247 1951 -213 1985
rect -247 1883 -213 1917
rect -247 1815 -213 1849
rect -247 1747 -213 1781
rect -247 1679 -213 1713
rect -247 1611 -213 1645
rect -247 1543 -213 1577
rect -247 1475 -213 1509
rect -247 1407 -213 1441
rect -247 1339 -213 1373
rect -247 1271 -213 1305
rect -247 1203 -213 1237
rect -247 1135 -213 1169
rect -247 1067 -213 1101
rect -247 999 -213 1033
rect -247 931 -213 965
rect -247 863 -213 897
rect -247 795 -213 829
rect -247 727 -213 761
rect -247 659 -213 693
rect -247 591 -213 625
rect -247 523 -213 557
rect -247 455 -213 489
rect -247 387 -213 421
rect -247 319 -213 353
rect -247 251 -213 285
rect -247 183 -213 217
rect -247 115 -213 149
rect -247 47 -213 81
rect -247 -21 -213 13
rect -247 -89 -213 -55
rect -247 -157 -213 -123
rect -247 -225 -213 -191
rect -247 -293 -213 -259
rect -247 -361 -213 -327
rect -247 -453 -213 -395
rect 4093 2835 4127 2883
rect 4093 2767 4127 2801
rect 4093 2699 4127 2733
rect 4093 2631 4127 2665
rect 4093 2563 4127 2597
rect 4093 2495 4127 2529
rect 4093 2427 4127 2461
rect 4093 2359 4127 2393
rect 4093 2291 4127 2325
rect 4093 2223 4127 2257
rect 4093 2155 4127 2189
rect 4093 2087 4127 2121
rect 4093 2019 4127 2053
rect 4093 1951 4127 1985
rect 4093 1883 4127 1917
rect 4093 1815 4127 1849
rect 4093 1747 4127 1781
rect 4093 1679 4127 1713
rect 4093 1611 4127 1645
rect 4093 1543 4127 1577
rect 4093 1475 4127 1509
rect 4093 1407 4127 1441
rect 4093 1339 4127 1373
rect 4093 1271 4127 1305
rect 4093 1203 4127 1237
rect 4093 1135 4127 1169
rect 4093 1067 4127 1101
rect 4093 999 4127 1033
rect 4093 931 4127 965
rect 4093 863 4127 897
rect 4093 795 4127 829
rect 4093 727 4127 761
rect 4093 659 4127 693
rect 4093 591 4127 625
rect 4093 523 4127 557
rect 4093 455 4127 489
rect 4093 387 4127 421
rect 4093 319 4127 353
rect 4093 251 4127 285
rect 4093 183 4127 217
rect 4093 115 4127 149
rect 4093 47 4127 81
rect 4093 -21 4127 13
rect 4093 -89 4127 -55
rect 4093 -157 4127 -123
rect 4093 -225 4127 -191
rect 4093 -293 4127 -259
rect 4093 -361 4127 -327
rect 4093 -453 4127 -395
rect -247 -487 -185 -453
rect -151 -487 -117 -453
rect -83 -487 -49 -453
rect -15 -487 19 -453
rect 53 -487 87 -453
rect 121 -487 155 -453
rect 189 -487 223 -453
rect 257 -487 291 -453
rect 325 -487 359 -453
rect 393 -487 427 -453
rect 461 -487 495 -453
rect 529 -487 563 -453
rect 597 -487 631 -453
rect 665 -487 699 -453
rect 733 -487 767 -453
rect 801 -487 835 -453
rect 869 -487 903 -453
rect 937 -487 971 -453
rect 1005 -487 1039 -453
rect 1073 -487 1107 -453
rect 1141 -487 1175 -453
rect 1209 -487 1243 -453
rect 1277 -487 1311 -453
rect 1345 -487 1379 -453
rect 1413 -487 1447 -453
rect 1481 -487 1515 -453
rect 1549 -487 1583 -453
rect 1617 -487 1651 -453
rect 1685 -487 1719 -453
rect 1753 -487 1787 -453
rect 1821 -487 1855 -453
rect 1889 -487 1923 -453
rect 1957 -487 1991 -453
rect 2025 -487 2059 -453
rect 2093 -487 2127 -453
rect 2161 -487 2195 -453
rect 2229 -487 2263 -453
rect 2297 -487 2331 -453
rect 2365 -487 2399 -453
rect 2433 -487 2467 -453
rect 2501 -487 2535 -453
rect 2569 -487 2603 -453
rect 2637 -487 2671 -453
rect 2705 -487 2739 -453
rect 2773 -487 2807 -453
rect 2841 -487 2875 -453
rect 2909 -487 2943 -453
rect 2977 -487 3011 -453
rect 3045 -487 3079 -453
rect 3113 -487 3147 -453
rect 3181 -487 3215 -453
rect 3249 -487 3283 -453
rect 3317 -487 3351 -453
rect 3385 -487 3419 -453
rect 3453 -487 3487 -453
rect 3521 -487 3555 -453
rect 3589 -487 3623 -453
rect 3657 -487 3691 -453
rect 3725 -487 3759 -453
rect 3793 -487 3827 -453
rect 3861 -487 3895 -453
rect 3929 -487 3963 -453
rect 3997 -487 4031 -453
rect 4065 -487 4127 -453
<< nsubdiffcont >>
rect -185 2883 -151 2917
rect -117 2883 -83 2917
rect -49 2883 -15 2917
rect 19 2883 53 2917
rect 87 2883 121 2917
rect 155 2883 189 2917
rect 223 2883 257 2917
rect 291 2883 325 2917
rect 359 2883 393 2917
rect 427 2883 461 2917
rect 495 2883 529 2917
rect 563 2883 597 2917
rect 631 2883 665 2917
rect 699 2883 733 2917
rect 767 2883 801 2917
rect 835 2883 869 2917
rect 903 2883 937 2917
rect 971 2883 1005 2917
rect 1039 2883 1073 2917
rect 1107 2883 1141 2917
rect 1175 2883 1209 2917
rect 1243 2883 1277 2917
rect 1311 2883 1345 2917
rect 1379 2883 1413 2917
rect 1447 2883 1481 2917
rect 1515 2883 1549 2917
rect 1583 2883 1617 2917
rect 1651 2883 1685 2917
rect 1719 2883 1753 2917
rect 1787 2883 1821 2917
rect 1855 2883 1889 2917
rect 1923 2883 1957 2917
rect 1991 2883 2025 2917
rect 2059 2883 2093 2917
rect 2127 2883 2161 2917
rect 2195 2883 2229 2917
rect 2263 2883 2297 2917
rect 2331 2883 2365 2917
rect 2399 2883 2433 2917
rect 2467 2883 2501 2917
rect 2535 2883 2569 2917
rect 2603 2883 2637 2917
rect 2671 2883 2705 2917
rect 2739 2883 2773 2917
rect 2807 2883 2841 2917
rect 2875 2883 2909 2917
rect 2943 2883 2977 2917
rect 3011 2883 3045 2917
rect 3079 2883 3113 2917
rect 3147 2883 3181 2917
rect 3215 2883 3249 2917
rect 3283 2883 3317 2917
rect 3351 2883 3385 2917
rect 3419 2883 3453 2917
rect 3487 2883 3521 2917
rect 3555 2883 3589 2917
rect 3623 2883 3657 2917
rect 3691 2883 3725 2917
rect 3759 2883 3793 2917
rect 3827 2883 3861 2917
rect 3895 2883 3929 2917
rect 3963 2883 3997 2917
rect 4031 2883 4065 2917
rect -247 2801 -213 2835
rect -247 2733 -213 2767
rect -247 2665 -213 2699
rect -247 2597 -213 2631
rect -247 2529 -213 2563
rect -247 2461 -213 2495
rect -247 2393 -213 2427
rect -247 2325 -213 2359
rect -247 2257 -213 2291
rect -247 2189 -213 2223
rect -247 2121 -213 2155
rect -247 2053 -213 2087
rect -247 1985 -213 2019
rect -247 1917 -213 1951
rect -247 1849 -213 1883
rect -247 1781 -213 1815
rect -247 1713 -213 1747
rect -247 1645 -213 1679
rect -247 1577 -213 1611
rect -247 1509 -213 1543
rect -247 1441 -213 1475
rect -247 1373 -213 1407
rect -247 1305 -213 1339
rect -247 1237 -213 1271
rect -247 1169 -213 1203
rect -247 1101 -213 1135
rect -247 1033 -213 1067
rect -247 965 -213 999
rect -247 897 -213 931
rect -247 829 -213 863
rect -247 761 -213 795
rect -247 693 -213 727
rect -247 625 -213 659
rect -247 557 -213 591
rect -247 489 -213 523
rect -247 421 -213 455
rect -247 353 -213 387
rect -247 285 -213 319
rect -247 217 -213 251
rect -247 149 -213 183
rect -247 81 -213 115
rect -247 13 -213 47
rect -247 -55 -213 -21
rect -247 -123 -213 -89
rect -247 -191 -213 -157
rect -247 -259 -213 -225
rect -247 -327 -213 -293
rect -247 -395 -213 -361
rect 4093 2801 4127 2835
rect 4093 2733 4127 2767
rect 4093 2665 4127 2699
rect 4093 2597 4127 2631
rect 4093 2529 4127 2563
rect 4093 2461 4127 2495
rect 4093 2393 4127 2427
rect 4093 2325 4127 2359
rect 4093 2257 4127 2291
rect 4093 2189 4127 2223
rect 4093 2121 4127 2155
rect 4093 2053 4127 2087
rect 4093 1985 4127 2019
rect 4093 1917 4127 1951
rect 4093 1849 4127 1883
rect 4093 1781 4127 1815
rect 4093 1713 4127 1747
rect 4093 1645 4127 1679
rect 4093 1577 4127 1611
rect 4093 1509 4127 1543
rect 4093 1441 4127 1475
rect 4093 1373 4127 1407
rect 4093 1305 4127 1339
rect 4093 1237 4127 1271
rect 4093 1169 4127 1203
rect 4093 1101 4127 1135
rect 4093 1033 4127 1067
rect 4093 965 4127 999
rect 4093 897 4127 931
rect 4093 829 4127 863
rect 4093 761 4127 795
rect 4093 693 4127 727
rect 4093 625 4127 659
rect 4093 557 4127 591
rect 4093 489 4127 523
rect 4093 421 4127 455
rect 4093 353 4127 387
rect 4093 285 4127 319
rect 4093 217 4127 251
rect 4093 149 4127 183
rect 4093 81 4127 115
rect 4093 13 4127 47
rect 4093 -55 4127 -21
rect 4093 -123 4127 -89
rect 4093 -191 4127 -157
rect 4093 -259 4127 -225
rect 4093 -327 4127 -293
rect 4093 -395 4127 -361
rect -185 -487 -151 -453
rect -117 -487 -83 -453
rect -49 -487 -15 -453
rect 19 -487 53 -453
rect 87 -487 121 -453
rect 155 -487 189 -453
rect 223 -487 257 -453
rect 291 -487 325 -453
rect 359 -487 393 -453
rect 427 -487 461 -453
rect 495 -487 529 -453
rect 563 -487 597 -453
rect 631 -487 665 -453
rect 699 -487 733 -453
rect 767 -487 801 -453
rect 835 -487 869 -453
rect 903 -487 937 -453
rect 971 -487 1005 -453
rect 1039 -487 1073 -453
rect 1107 -487 1141 -453
rect 1175 -487 1209 -453
rect 1243 -487 1277 -453
rect 1311 -487 1345 -453
rect 1379 -487 1413 -453
rect 1447 -487 1481 -453
rect 1515 -487 1549 -453
rect 1583 -487 1617 -453
rect 1651 -487 1685 -453
rect 1719 -487 1753 -453
rect 1787 -487 1821 -453
rect 1855 -487 1889 -453
rect 1923 -487 1957 -453
rect 1991 -487 2025 -453
rect 2059 -487 2093 -453
rect 2127 -487 2161 -453
rect 2195 -487 2229 -453
rect 2263 -487 2297 -453
rect 2331 -487 2365 -453
rect 2399 -487 2433 -453
rect 2467 -487 2501 -453
rect 2535 -487 2569 -453
rect 2603 -487 2637 -453
rect 2671 -487 2705 -453
rect 2739 -487 2773 -453
rect 2807 -487 2841 -453
rect 2875 -487 2909 -453
rect 2943 -487 2977 -453
rect 3011 -487 3045 -453
rect 3079 -487 3113 -453
rect 3147 -487 3181 -453
rect 3215 -487 3249 -453
rect 3283 -487 3317 -453
rect 3351 -487 3385 -453
rect 3419 -487 3453 -453
rect 3487 -487 3521 -453
rect 3555 -487 3589 -453
rect 3623 -487 3657 -453
rect 3691 -487 3725 -453
rect 3759 -487 3793 -453
rect 3827 -487 3861 -453
rect 3895 -487 3929 -453
rect 3963 -487 3997 -453
rect 4031 -487 4065 -453
<< locali >>
rect -247 2883 -185 2917
rect -151 2883 -117 2917
rect -83 2883 -49 2917
rect -15 2883 19 2917
rect 53 2883 87 2917
rect 121 2883 155 2917
rect 189 2883 223 2917
rect 257 2883 291 2917
rect 325 2883 359 2917
rect 393 2883 427 2917
rect 461 2883 495 2917
rect 529 2883 563 2917
rect 597 2883 631 2917
rect 665 2883 699 2917
rect 733 2883 767 2917
rect 801 2883 835 2917
rect 869 2883 903 2917
rect 937 2883 971 2917
rect 1005 2883 1039 2917
rect 1073 2883 1107 2917
rect 1141 2883 1175 2917
rect 1209 2883 1243 2917
rect 1277 2883 1311 2917
rect 1345 2883 1379 2917
rect 1413 2883 1447 2917
rect 1481 2883 1515 2917
rect 1549 2883 1583 2917
rect 1617 2883 1651 2917
rect 1685 2883 1719 2917
rect 1753 2883 1787 2917
rect 1821 2883 1855 2917
rect 1889 2883 1923 2917
rect 1957 2883 1991 2917
rect 2025 2883 2059 2917
rect 2093 2883 2127 2917
rect 2161 2883 2195 2917
rect 2229 2883 2263 2917
rect 2297 2883 2331 2917
rect 2365 2883 2399 2917
rect 2433 2883 2467 2917
rect 2501 2883 2535 2917
rect 2569 2883 2603 2917
rect 2637 2883 2671 2917
rect 2705 2883 2739 2917
rect 2773 2883 2807 2917
rect 2841 2883 2875 2917
rect 2909 2883 2943 2917
rect 2977 2883 3011 2917
rect 3045 2883 3079 2917
rect 3113 2883 3147 2917
rect 3181 2883 3215 2917
rect 3249 2883 3283 2917
rect 3317 2883 3351 2917
rect 3385 2883 3419 2917
rect 3453 2883 3487 2917
rect 3521 2883 3555 2917
rect 3589 2883 3623 2917
rect 3657 2883 3691 2917
rect 3725 2883 3759 2917
rect 3793 2883 3827 2917
rect 3861 2883 3895 2917
rect 3929 2883 3963 2917
rect 3997 2883 4031 2917
rect 4065 2883 4127 2917
rect -247 2835 -213 2883
rect -247 2767 -213 2801
rect -247 2699 -213 2733
rect -247 2631 -213 2665
rect -247 2563 -213 2597
rect -247 2495 -213 2529
rect -247 2427 -213 2461
rect -247 2359 -213 2393
rect -247 2291 -213 2325
rect -247 2223 -213 2257
rect -247 2155 -213 2189
rect -247 2087 -213 2121
rect -247 2019 -213 2053
rect -247 1951 -213 1985
rect -247 1883 -213 1917
rect -247 1815 -213 1849
rect -247 1747 -213 1781
rect -247 1679 -213 1713
rect -247 1611 -213 1645
rect -247 1543 -213 1577
rect -247 1475 -213 1509
rect -247 1407 -213 1441
rect -247 1339 -213 1373
rect -247 1271 -213 1305
rect -247 1203 -213 1237
rect -247 1135 -213 1169
rect -247 1067 -213 1101
rect -247 999 -213 1033
rect -247 931 -213 965
rect -247 863 -213 897
rect -247 795 -213 829
rect -247 727 -213 761
rect -247 659 -213 693
rect -247 591 -213 625
rect -247 523 -213 557
rect -247 455 -213 489
rect -247 387 -213 421
rect -247 319 -213 353
rect -247 251 -213 285
rect -247 183 -213 217
rect -247 115 -213 149
rect -247 47 -213 81
rect -247 -21 -213 13
rect -247 -89 -213 -55
rect -247 -157 -213 -123
rect -247 -225 -213 -191
rect -247 -293 -213 -259
rect -247 -361 -213 -327
rect -247 -453 -213 -395
rect 4093 2835 4127 2883
rect 4093 2767 4127 2801
rect 4093 2699 4127 2733
rect 4093 2631 4127 2665
rect 4093 2563 4127 2597
rect 4093 2495 4127 2529
rect 4093 2427 4127 2461
rect 4093 2359 4127 2393
rect 4093 2291 4127 2325
rect 4093 2223 4127 2257
rect 4093 2155 4127 2189
rect 4093 2087 4127 2121
rect 4093 2019 4127 2053
rect 4093 1951 4127 1985
rect 4093 1883 4127 1917
rect 4093 1815 4127 1849
rect 4093 1747 4127 1781
rect 4093 1679 4127 1713
rect 4093 1611 4127 1645
rect 4093 1543 4127 1577
rect 4093 1475 4127 1509
rect 4093 1407 4127 1441
rect 4093 1339 4127 1373
rect 4093 1271 4127 1305
rect 4093 1203 4127 1237
rect 4093 1135 4127 1169
rect 4093 1067 4127 1101
rect 4093 999 4127 1033
rect 4093 931 4127 965
rect 4093 863 4127 897
rect 4093 795 4127 829
rect 4093 727 4127 761
rect 4093 659 4127 693
rect 4093 591 4127 625
rect 4093 523 4127 557
rect 4093 455 4127 489
rect 4093 387 4127 421
rect 4093 319 4127 353
rect 4093 251 4127 285
rect 4093 183 4127 217
rect 4093 115 4127 149
rect 4093 47 4127 81
rect 4093 -21 4127 13
rect 4093 -89 4127 -55
rect 4093 -157 4127 -123
rect 4093 -225 4127 -191
rect 4093 -293 4127 -259
rect 4093 -361 4127 -327
rect 4093 -453 4127 -395
rect -247 -487 -185 -453
rect -151 -487 -117 -453
rect -83 -487 -49 -453
rect -15 -487 19 -453
rect 53 -487 87 -453
rect 121 -487 155 -453
rect 189 -487 223 -453
rect 257 -487 291 -453
rect 325 -487 359 -453
rect 393 -487 427 -453
rect 461 -487 495 -453
rect 529 -487 563 -453
rect 597 -487 631 -453
rect 665 -487 699 -453
rect 733 -487 767 -453
rect 801 -487 835 -453
rect 869 -487 903 -453
rect 937 -487 971 -453
rect 1005 -487 1039 -453
rect 1073 -487 1107 -453
rect 1141 -487 1175 -453
rect 1209 -487 1243 -453
rect 1277 -487 1311 -453
rect 1345 -487 1379 -453
rect 1413 -487 1447 -453
rect 1481 -487 1515 -453
rect 1549 -487 1583 -453
rect 1617 -487 1651 -453
rect 1685 -487 1719 -453
rect 1753 -487 1787 -453
rect 1821 -487 1855 -453
rect 1889 -487 1923 -453
rect 1957 -487 1991 -453
rect 2025 -487 2059 -453
rect 2093 -487 2127 -453
rect 2161 -487 2195 -453
rect 2229 -487 2263 -453
rect 2297 -487 2331 -453
rect 2365 -487 2399 -453
rect 2433 -487 2467 -453
rect 2501 -487 2535 -453
rect 2569 -487 2603 -453
rect 2637 -487 2671 -453
rect 2705 -487 2739 -453
rect 2773 -487 2807 -453
rect 2841 -487 2875 -453
rect 2909 -487 2943 -453
rect 2977 -487 3011 -453
rect 3045 -487 3079 -453
rect 3113 -487 3147 -453
rect 3181 -487 3215 -453
rect 3249 -487 3283 -453
rect 3317 -487 3351 -453
rect 3385 -487 3419 -453
rect 3453 -487 3487 -453
rect 3521 -487 3555 -453
rect 3589 -487 3623 -453
rect 3657 -487 3691 -453
rect 3725 -487 3759 -453
rect 3793 -487 3827 -453
rect 3861 -487 3895 -453
rect 3929 -487 3963 -453
rect 3997 -487 4031 -453
rect 4065 -487 4127 -453
<< metal1 >>
rect 60 3020 280 3030
rect 60 2710 3950 3020
rect 280 2520 3950 2710
rect 60 2460 3950 2520
rect 60 2380 250 2460
rect 3680 2380 3950 2460
rect 60 2376 350 2380
rect 60 2324 89 2376
rect 141 2324 350 2376
rect 60 2320 350 2324
rect 460 2376 660 2380
rect 460 2324 484 2376
rect 536 2324 584 2376
rect 636 2324 660 2376
rect 460 2320 660 2324
rect 860 2376 1060 2380
rect 860 2324 884 2376
rect 936 2324 984 2376
rect 1036 2324 1060 2376
rect 860 2320 1060 2324
rect 1260 2376 1460 2380
rect 1260 2324 1284 2376
rect 1336 2324 1384 2376
rect 1436 2324 1460 2376
rect 1260 2320 1460 2324
rect 1660 2376 1860 2380
rect 1660 2324 1684 2376
rect 1736 2324 1784 2376
rect 1836 2324 1860 2376
rect 1660 2320 1860 2324
rect 2060 2376 2260 2380
rect 2060 2324 2084 2376
rect 2136 2324 2184 2376
rect 2236 2324 2260 2376
rect 2060 2320 2260 2324
rect 2460 2376 2660 2380
rect 2460 2324 2484 2376
rect 2536 2324 2584 2376
rect 2636 2324 2660 2376
rect 2460 2320 2660 2324
rect 2860 2376 3060 2380
rect 2860 2324 2884 2376
rect 2936 2324 2984 2376
rect 3036 2324 3060 2376
rect 2860 2320 3060 2324
rect 3260 2376 3460 2380
rect 3260 2324 3284 2376
rect 3336 2324 3384 2376
rect 3436 2324 3460 2376
rect 3260 2320 3460 2324
rect 3660 2376 3950 2380
rect 3660 2324 3694 2376
rect 3746 2324 3794 2376
rect 3846 2324 3950 2376
rect 3660 2320 3950 2324
rect -60 1406 20 1410
rect -60 1354 -46 1406
rect 6 1354 20 1406
rect -60 1326 20 1354
rect 290 1330 350 2320
rect 670 2016 750 2040
rect 670 1964 684 2016
rect 736 1964 750 2016
rect 670 1926 750 1964
rect 670 1874 684 1926
rect 736 1874 750 1926
rect 670 1836 750 1874
rect 670 1784 684 1836
rect 736 1784 750 1836
rect 670 1746 750 1784
rect 670 1694 684 1746
rect 736 1694 750 1746
rect 670 1680 750 1694
rect 1070 2016 1150 2040
rect 1070 1964 1084 2016
rect 1136 1964 1150 2016
rect 1070 1926 1150 1964
rect 1070 1874 1084 1926
rect 1136 1874 1150 1926
rect 1070 1836 1150 1874
rect 1070 1784 1084 1836
rect 1136 1784 1150 1836
rect 1070 1746 1150 1784
rect 1070 1694 1084 1746
rect 1136 1694 1150 1746
rect 1070 1680 1150 1694
rect 1470 2016 1550 2040
rect 1470 1964 1484 2016
rect 1536 1964 1550 2016
rect 1470 1926 1550 1964
rect 1470 1874 1484 1926
rect 1536 1874 1550 1926
rect 1470 1836 1550 1874
rect 1470 1784 1484 1836
rect 1536 1784 1550 1836
rect 1470 1746 1550 1784
rect 1470 1694 1484 1746
rect 1536 1694 1550 1746
rect 1470 1680 1550 1694
rect 1870 2016 1950 2040
rect 1870 1964 1884 2016
rect 1936 1964 1950 2016
rect 1870 1926 1950 1964
rect 1870 1874 1884 1926
rect 1936 1874 1950 1926
rect 1870 1836 1950 1874
rect 1870 1784 1884 1836
rect 1936 1784 1950 1836
rect 1870 1746 1950 1784
rect 1870 1694 1884 1746
rect 1936 1694 1950 1746
rect 1870 1680 1950 1694
rect 2270 2016 2350 2040
rect 2270 1964 2284 2016
rect 2336 1964 2350 2016
rect 2270 1926 2350 1964
rect 2270 1874 2284 1926
rect 2336 1874 2350 1926
rect 2270 1836 2350 1874
rect 2270 1784 2284 1836
rect 2336 1784 2350 1836
rect 2270 1746 2350 1784
rect 2270 1694 2284 1746
rect 2336 1694 2350 1746
rect 2270 1680 2350 1694
rect 2670 2016 2750 2040
rect 2670 1964 2684 2016
rect 2736 1964 2750 2016
rect 2670 1926 2750 1964
rect 2670 1874 2684 1926
rect 2736 1874 2750 1926
rect 2670 1836 2750 1874
rect 2670 1784 2684 1836
rect 2736 1784 2750 1836
rect 2670 1746 2750 1784
rect 2670 1694 2684 1746
rect 2736 1694 2750 1746
rect 2670 1680 2750 1694
rect 3070 2016 3150 2040
rect 3070 1964 3084 2016
rect 3136 1964 3150 2016
rect 3070 1926 3150 1964
rect 3070 1874 3084 1926
rect 3136 1874 3150 1926
rect 3070 1836 3150 1874
rect 3070 1784 3084 1836
rect 3136 1784 3150 1836
rect 3070 1746 3150 1784
rect 3070 1694 3084 1746
rect 3136 1694 3150 1746
rect 3070 1680 3150 1694
rect 3470 2016 3550 2040
rect 3470 1964 3484 2016
rect 3536 1964 3550 2016
rect 3470 1926 3550 1964
rect 3470 1874 3484 1926
rect 3536 1874 3550 1926
rect 3470 1836 3550 1874
rect 3470 1784 3484 1836
rect 3536 1784 3550 1836
rect 3470 1746 3550 1784
rect 3470 1694 3484 1746
rect 3536 1694 3550 1746
rect 3470 1680 3550 1694
rect 3890 1330 3950 2320
rect -60 1274 -46 1326
rect 6 1274 20 1326
rect -60 176 20 1274
rect 60 1146 350 1330
rect 470 1326 650 1330
rect 470 1274 494 1326
rect 546 1274 574 1326
rect 626 1274 650 1326
rect 470 1270 650 1274
rect 870 1326 1050 1330
rect 870 1274 894 1326
rect 946 1274 974 1326
rect 1026 1274 1050 1326
rect 870 1270 1050 1274
rect 1270 1236 1450 1330
rect 1270 1184 1294 1236
rect 1346 1184 1374 1236
rect 1426 1184 1450 1236
rect 1270 1180 1450 1184
rect 1670 1236 1850 1330
rect 1670 1184 1694 1236
rect 1746 1184 1774 1236
rect 1826 1184 1850 1236
rect 1670 1180 1850 1184
rect 2070 1236 2250 1330
rect 2070 1184 2094 1236
rect 2146 1184 2174 1236
rect 2226 1184 2250 1236
rect 2070 1180 2250 1184
rect 2470 1236 2650 1330
rect 2870 1326 3050 1330
rect 2870 1274 2894 1326
rect 2946 1274 2974 1326
rect 3026 1274 3050 1326
rect 2870 1270 3050 1274
rect 3270 1326 3450 1330
rect 3270 1274 3294 1326
rect 3346 1274 3374 1326
rect 3426 1274 3450 1326
rect 3270 1270 3450 1274
rect 2470 1184 2494 1236
rect 2546 1184 2574 1236
rect 2626 1184 2650 1236
rect 2470 1180 2650 1184
rect 60 1094 94 1146
rect 146 1094 194 1146
rect 246 1094 350 1146
rect 60 1090 350 1094
rect 470 1146 650 1150
rect 470 1094 484 1146
rect 536 1094 574 1146
rect 626 1094 650 1146
rect 470 1090 650 1094
rect 870 1146 1050 1150
rect 870 1094 894 1146
rect 946 1094 974 1146
rect 1026 1094 1050 1146
rect 870 1090 1050 1094
rect 1270 1146 1450 1150
rect 1270 1094 1294 1146
rect 1346 1094 1374 1146
rect 1426 1094 1450 1146
rect 1270 1090 1450 1094
rect 1670 1146 1850 1150
rect 1670 1094 1694 1146
rect 1746 1094 1774 1146
rect 1826 1094 1850 1146
rect 1670 1090 1850 1094
rect 2070 1146 2250 1150
rect 2070 1094 2094 1146
rect 2146 1094 2174 1146
rect 2226 1094 2250 1146
rect 2070 1090 2250 1094
rect 2470 1146 2650 1150
rect 2470 1094 2494 1146
rect 2546 1094 2574 1146
rect 2626 1094 2650 1146
rect 2470 1090 2650 1094
rect 2870 1146 3050 1150
rect 2870 1094 2894 1146
rect 2946 1094 2974 1146
rect 3026 1094 3050 1146
rect 2870 1090 3050 1094
rect 3270 1146 3450 1150
rect 3270 1094 3294 1146
rect 3346 1094 3374 1146
rect 3426 1094 3450 1146
rect 3270 1090 3450 1094
rect 3660 1146 3950 1330
rect 3660 1094 3684 1146
rect 3736 1094 3774 1146
rect 3826 1094 3950 1146
rect 3660 1090 3950 1094
rect -60 124 -46 176
rect 6 124 20 176
rect -60 96 20 124
rect 290 100 350 1090
rect 670 796 750 820
rect 670 744 684 796
rect 736 744 750 796
rect 670 706 750 744
rect 670 654 684 706
rect 736 654 750 706
rect 670 616 750 654
rect 670 564 684 616
rect 736 564 750 616
rect 670 526 750 564
rect 670 474 684 526
rect 736 474 750 526
rect 670 460 750 474
rect 1070 796 1150 820
rect 1070 744 1084 796
rect 1136 744 1150 796
rect 1070 706 1150 744
rect 1070 654 1084 706
rect 1136 654 1150 706
rect 1070 616 1150 654
rect 1070 564 1084 616
rect 1136 564 1150 616
rect 1070 526 1150 564
rect 1070 474 1084 526
rect 1136 474 1150 526
rect 1070 460 1150 474
rect 1470 796 1550 820
rect 1470 744 1484 796
rect 1536 744 1550 796
rect 1470 706 1550 744
rect 1470 654 1484 706
rect 1536 654 1550 706
rect 1470 616 1550 654
rect 1470 564 1484 616
rect 1536 564 1550 616
rect 1470 526 1550 564
rect 1470 474 1484 526
rect 1536 474 1550 526
rect 1470 460 1550 474
rect 1870 796 1950 820
rect 1870 744 1884 796
rect 1936 744 1950 796
rect 1870 706 1950 744
rect 1870 654 1884 706
rect 1936 654 1950 706
rect 1870 616 1950 654
rect 1870 564 1884 616
rect 1936 564 1950 616
rect 1870 526 1950 564
rect 1870 474 1884 526
rect 1936 474 1950 526
rect 1870 460 1950 474
rect 2270 796 2350 820
rect 2270 744 2284 796
rect 2336 744 2350 796
rect 2270 706 2350 744
rect 2270 654 2284 706
rect 2336 654 2350 706
rect 2270 616 2350 654
rect 2270 564 2284 616
rect 2336 564 2350 616
rect 2270 526 2350 564
rect 2270 474 2284 526
rect 2336 474 2350 526
rect 2270 460 2350 474
rect 2670 796 2750 820
rect 2670 744 2684 796
rect 2736 744 2750 796
rect 2670 706 2750 744
rect 2670 654 2684 706
rect 2736 654 2750 706
rect 2670 616 2750 654
rect 2670 564 2684 616
rect 2736 564 2750 616
rect 2670 526 2750 564
rect 2670 474 2684 526
rect 2736 474 2750 526
rect 2670 460 2750 474
rect 3070 796 3150 820
rect 3070 744 3084 796
rect 3136 744 3150 796
rect 3070 706 3150 744
rect 3070 654 3084 706
rect 3136 654 3150 706
rect 3070 616 3150 654
rect 3070 564 3084 616
rect 3136 564 3150 616
rect 3070 526 3150 564
rect 3070 474 3084 526
rect 3136 474 3150 526
rect 3070 460 3150 474
rect 3470 796 3550 820
rect 3470 744 3484 796
rect 3536 744 3550 796
rect 3470 706 3550 744
rect 3470 654 3484 706
rect 3536 654 3550 706
rect 3470 616 3550 654
rect 3470 564 3484 616
rect 3536 564 3550 616
rect 3470 526 3550 564
rect 3470 474 3484 526
rect 3536 474 3550 526
rect 3470 460 3550 474
rect 3890 100 3950 1090
rect -60 44 -46 96
rect 6 44 20 96
rect -60 40 20 44
rect 60 -80 350 100
rect 470 6 650 100
rect 470 -46 494 6
rect 546 -46 574 6
rect 626 -46 650 6
rect 470 -50 650 -46
rect 870 6 1050 100
rect 1270 96 1450 100
rect 1270 44 1294 96
rect 1346 44 1374 96
rect 1426 44 1450 96
rect 1270 40 1450 44
rect 1670 96 1850 100
rect 1670 44 1694 96
rect 1746 44 1774 96
rect 1826 44 1850 96
rect 1670 40 1850 44
rect 2070 96 2250 100
rect 2070 44 2094 96
rect 2146 44 2174 96
rect 2226 44 2250 96
rect 2070 40 2250 44
rect 2470 96 2650 100
rect 2470 44 2494 96
rect 2546 44 2574 96
rect 2626 44 2650 96
rect 2470 40 2650 44
rect 870 -46 894 6
rect 946 -46 974 6
rect 1026 -46 1050 6
rect 870 -50 1050 -46
rect 2870 6 3050 100
rect 2870 -46 2894 6
rect 2946 -46 2974 6
rect 3026 -46 3050 6
rect 2870 -50 3050 -46
rect 3270 6 3450 100
rect 3270 -46 3294 6
rect 3346 -46 3374 6
rect 3426 -46 3450 6
rect 3270 -50 3450 -46
rect 3660 -80 3950 100
rect 3980 1236 4060 1240
rect 3980 1184 3994 1236
rect 4046 1184 4060 1236
rect 3980 1156 4060 1184
rect 3980 1104 3994 1156
rect 4046 1104 4060 1156
rect 3980 86 4060 1104
rect 3980 34 3994 86
rect 4046 34 4060 86
rect 3980 6 4060 34
rect 3980 -46 3994 6
rect 4046 -46 4060 6
rect 3980 -50 4060 -46
rect 60 -390 3950 -80
<< via1 >>
rect 89 2324 141 2376
rect 484 2324 536 2376
rect 584 2324 636 2376
rect 884 2324 936 2376
rect 984 2324 1036 2376
rect 1284 2324 1336 2376
rect 1384 2324 1436 2376
rect 1684 2324 1736 2376
rect 1784 2324 1836 2376
rect 2084 2324 2136 2376
rect 2184 2324 2236 2376
rect 2484 2324 2536 2376
rect 2584 2324 2636 2376
rect 2884 2324 2936 2376
rect 2984 2324 3036 2376
rect 3284 2324 3336 2376
rect 3384 2324 3436 2376
rect 3694 2324 3746 2376
rect 3794 2324 3846 2376
rect -46 1354 6 1406
rect 684 1964 736 2016
rect 684 1874 736 1926
rect 684 1784 736 1836
rect 684 1694 736 1746
rect 1084 1964 1136 2016
rect 1084 1874 1136 1926
rect 1084 1784 1136 1836
rect 1084 1694 1136 1746
rect 1484 1964 1536 2016
rect 1484 1874 1536 1926
rect 1484 1784 1536 1836
rect 1484 1694 1536 1746
rect 1884 1964 1936 2016
rect 1884 1874 1936 1926
rect 1884 1784 1936 1836
rect 1884 1694 1936 1746
rect 2284 1964 2336 2016
rect 2284 1874 2336 1926
rect 2284 1784 2336 1836
rect 2284 1694 2336 1746
rect 2684 1964 2736 2016
rect 2684 1874 2736 1926
rect 2684 1784 2736 1836
rect 2684 1694 2736 1746
rect 3084 1964 3136 2016
rect 3084 1874 3136 1926
rect 3084 1784 3136 1836
rect 3084 1694 3136 1746
rect 3484 1964 3536 2016
rect 3484 1874 3536 1926
rect 3484 1784 3536 1836
rect 3484 1694 3536 1746
rect -46 1274 6 1326
rect 494 1274 546 1326
rect 574 1274 626 1326
rect 894 1274 946 1326
rect 974 1274 1026 1326
rect 1294 1184 1346 1236
rect 1374 1184 1426 1236
rect 1694 1184 1746 1236
rect 1774 1184 1826 1236
rect 2094 1184 2146 1236
rect 2174 1184 2226 1236
rect 2894 1274 2946 1326
rect 2974 1274 3026 1326
rect 3294 1274 3346 1326
rect 3374 1274 3426 1326
rect 2494 1184 2546 1236
rect 2574 1184 2626 1236
rect 94 1094 146 1146
rect 194 1094 246 1146
rect 484 1094 536 1146
rect 574 1094 626 1146
rect 894 1094 946 1146
rect 974 1094 1026 1146
rect 1294 1094 1346 1146
rect 1374 1094 1426 1146
rect 1694 1094 1746 1146
rect 1774 1094 1826 1146
rect 2094 1094 2146 1146
rect 2174 1094 2226 1146
rect 2494 1094 2546 1146
rect 2574 1094 2626 1146
rect 2894 1094 2946 1146
rect 2974 1094 3026 1146
rect 3294 1094 3346 1146
rect 3374 1094 3426 1146
rect 3684 1094 3736 1146
rect 3774 1094 3826 1146
rect -46 124 6 176
rect 684 744 736 796
rect 684 654 736 706
rect 684 564 736 616
rect 684 474 736 526
rect 1084 744 1136 796
rect 1084 654 1136 706
rect 1084 564 1136 616
rect 1084 474 1136 526
rect 1484 744 1536 796
rect 1484 654 1536 706
rect 1484 564 1536 616
rect 1484 474 1536 526
rect 1884 744 1936 796
rect 1884 654 1936 706
rect 1884 564 1936 616
rect 1884 474 1936 526
rect 2284 744 2336 796
rect 2284 654 2336 706
rect 2284 564 2336 616
rect 2284 474 2336 526
rect 2684 744 2736 796
rect 2684 654 2736 706
rect 2684 564 2736 616
rect 2684 474 2736 526
rect 3084 744 3136 796
rect 3084 654 3136 706
rect 3084 564 3136 616
rect 3084 474 3136 526
rect 3484 744 3536 796
rect 3484 654 3536 706
rect 3484 564 3536 616
rect 3484 474 3536 526
rect -46 44 6 96
rect 494 -46 546 6
rect 574 -46 626 6
rect 1294 44 1346 96
rect 1374 44 1426 96
rect 1694 44 1746 96
rect 1774 44 1826 96
rect 2094 44 2146 96
rect 2174 44 2226 96
rect 2494 44 2546 96
rect 2574 44 2626 96
rect 894 -46 946 6
rect 974 -46 1026 6
rect 2894 -46 2946 6
rect 2974 -46 3026 6
rect 3294 -46 3346 6
rect 3374 -46 3426 6
rect 3994 1184 4046 1236
rect 3994 1104 4046 1156
rect 3994 34 4046 86
rect 3994 -46 4046 6
<< metal2 >>
rect -80 2998 20 3020
rect -80 2942 -58 2998
rect -2 2942 20 2998
rect -80 2920 20 2942
rect -60 1406 20 2920
rect 4160 2860 4260 2870
rect 690 2848 4260 2860
rect 690 2792 702 2848
rect 758 2792 792 2848
rect 848 2792 1052 2848
rect 1108 2792 1142 2848
rect 1198 2792 1452 2848
rect 1508 2792 1542 2848
rect 1598 2792 1852 2848
rect 1908 2792 1942 2848
rect 1998 2792 2252 2848
rect 2308 2792 2342 2848
rect 2398 2792 2652 2848
rect 2708 2792 2742 2848
rect 2798 2792 3052 2848
rect 3108 2792 3142 2848
rect 3198 2792 3452 2848
rect 3508 2792 3542 2848
rect 3598 2792 4182 2848
rect 4238 2792 4260 2848
rect 690 2780 4260 2792
rect 4160 2770 4260 2780
rect 60 2376 3860 2380
rect 60 2324 89 2376
rect 141 2324 484 2376
rect 536 2324 584 2376
rect 636 2324 884 2376
rect 936 2324 984 2376
rect 1036 2324 1284 2376
rect 1336 2324 1384 2376
rect 1436 2324 1684 2376
rect 1736 2324 1784 2376
rect 1836 2324 2084 2376
rect 2136 2324 2184 2376
rect 2236 2324 2484 2376
rect 2536 2324 2584 2376
rect 2636 2324 2884 2376
rect 2936 2324 2984 2376
rect 3036 2324 3284 2376
rect 3336 2324 3384 2376
rect 3436 2324 3694 2376
rect 3746 2324 3794 2376
rect 3846 2324 3860 2376
rect 60 2320 3860 2324
rect 670 2018 750 2040
rect 670 1962 682 2018
rect 738 1962 750 2018
rect 670 1928 750 1962
rect 670 1872 682 1928
rect 738 1872 750 1928
rect 670 1838 750 1872
rect 670 1782 682 1838
rect 738 1782 750 1838
rect 670 1748 750 1782
rect 670 1692 682 1748
rect 738 1692 750 1748
rect 670 1680 750 1692
rect 1070 2018 1150 2040
rect 1070 1962 1082 2018
rect 1138 1962 1150 2018
rect 1070 1928 1150 1962
rect 1070 1872 1082 1928
rect 1138 1872 1150 1928
rect 1070 1838 1150 1872
rect 1070 1782 1082 1838
rect 1138 1782 1150 1838
rect 1070 1748 1150 1782
rect 1070 1692 1082 1748
rect 1138 1692 1150 1748
rect 1070 1680 1150 1692
rect 1470 2018 1550 2040
rect 1470 1962 1482 2018
rect 1538 1962 1550 2018
rect 1470 1928 1550 1962
rect 1470 1872 1482 1928
rect 1538 1872 1550 1928
rect 1470 1838 1550 1872
rect 1470 1782 1482 1838
rect 1538 1782 1550 1838
rect 1470 1748 1550 1782
rect 1470 1692 1482 1748
rect 1538 1692 1550 1748
rect 1470 1680 1550 1692
rect 1870 2018 1950 2040
rect 1870 1962 1882 2018
rect 1938 1962 1950 2018
rect 1870 1928 1950 1962
rect 1870 1872 1882 1928
rect 1938 1872 1950 1928
rect 1870 1838 1950 1872
rect 1870 1782 1882 1838
rect 1938 1782 1950 1838
rect 1870 1748 1950 1782
rect 1870 1692 1882 1748
rect 1938 1692 1950 1748
rect 1870 1680 1950 1692
rect 2270 2018 2350 2040
rect 2270 1962 2282 2018
rect 2338 1962 2350 2018
rect 2270 1928 2350 1962
rect 2270 1872 2282 1928
rect 2338 1872 2350 1928
rect 2270 1838 2350 1872
rect 2270 1782 2282 1838
rect 2338 1782 2350 1838
rect 2270 1748 2350 1782
rect 2270 1692 2282 1748
rect 2338 1692 2350 1748
rect 2270 1680 2350 1692
rect 2670 2018 2750 2040
rect 2670 1962 2682 2018
rect 2738 1962 2750 2018
rect 2670 1928 2750 1962
rect 2670 1872 2682 1928
rect 2738 1872 2750 1928
rect 2670 1838 2750 1872
rect 2670 1782 2682 1838
rect 2738 1782 2750 1838
rect 2670 1748 2750 1782
rect 2670 1692 2682 1748
rect 2738 1692 2750 1748
rect 2670 1680 2750 1692
rect 3070 2018 3150 2040
rect 3070 1962 3082 2018
rect 3138 1962 3150 2018
rect 3070 1928 3150 1962
rect 3070 1872 3082 1928
rect 3138 1872 3150 1928
rect 3070 1838 3150 1872
rect 3070 1782 3082 1838
rect 3138 1782 3150 1838
rect 3070 1748 3150 1782
rect 3070 1692 3082 1748
rect 3138 1692 3150 1748
rect 3070 1680 3150 1692
rect 3470 2018 3550 2040
rect 3470 1962 3482 2018
rect 3538 1962 3550 2018
rect 3470 1928 3550 1962
rect 3470 1872 3482 1928
rect 3538 1872 3550 1928
rect 3470 1838 3550 1872
rect 3470 1782 3482 1838
rect 3538 1782 3550 1838
rect 3470 1748 3550 1782
rect 3470 1692 3482 1748
rect 3538 1692 3550 1748
rect 3470 1680 3550 1692
rect -60 1354 -46 1406
rect 6 1354 20 1406
rect -60 1330 20 1354
rect -60 1326 3840 1330
rect -60 1274 -46 1326
rect 6 1274 494 1326
rect 546 1274 574 1326
rect 626 1274 894 1326
rect 946 1274 974 1326
rect 1026 1274 2894 1326
rect 2946 1274 2974 1326
rect 3026 1274 3294 1326
rect 3346 1274 3374 1326
rect 3426 1274 3840 1326
rect -60 1270 3840 1274
rect -180 1248 -100 1260
rect -180 1192 -168 1248
rect -112 1240 -100 1248
rect -112 1236 4060 1240
rect -112 1192 1294 1236
rect -180 1184 1294 1192
rect 1346 1184 1374 1236
rect 1426 1184 1694 1236
rect 1746 1184 1774 1236
rect 1826 1184 2094 1236
rect 2146 1184 2174 1236
rect 2226 1184 2494 1236
rect 2546 1184 2574 1236
rect 2626 1184 3994 1236
rect 4046 1184 4060 1236
rect -180 1180 4060 1184
rect 3980 1156 4060 1180
rect 60 1146 3840 1150
rect 60 1094 94 1146
rect 146 1094 194 1146
rect 246 1094 484 1146
rect 536 1094 574 1146
rect 626 1094 894 1146
rect 946 1094 974 1146
rect 1026 1094 1294 1146
rect 1346 1094 1374 1146
rect 1426 1094 1694 1146
rect 1746 1094 1774 1146
rect 1826 1094 2094 1146
rect 2146 1094 2174 1146
rect 2226 1094 2494 1146
rect 2546 1094 2574 1146
rect 2626 1094 2894 1146
rect 2946 1094 2974 1146
rect 3026 1094 3294 1146
rect 3346 1094 3374 1146
rect 3426 1094 3684 1146
rect 3736 1094 3774 1146
rect 3826 1094 3840 1146
rect 3980 1104 3994 1156
rect 4046 1104 4060 1156
rect 3980 1100 4060 1104
rect 60 1090 3840 1094
rect 670 798 750 820
rect 670 742 682 798
rect 738 742 750 798
rect 670 708 750 742
rect 670 652 682 708
rect 738 652 750 708
rect 670 618 750 652
rect 670 562 682 618
rect 738 562 750 618
rect 670 528 750 562
rect 670 472 682 528
rect 738 472 750 528
rect 670 460 750 472
rect 1070 798 1150 820
rect 1070 742 1082 798
rect 1138 742 1150 798
rect 1070 708 1150 742
rect 1070 652 1082 708
rect 1138 652 1150 708
rect 1070 618 1150 652
rect 1070 562 1082 618
rect 1138 562 1150 618
rect 1070 528 1150 562
rect 1070 472 1082 528
rect 1138 472 1150 528
rect 1070 460 1150 472
rect 1470 798 1550 820
rect 1470 742 1482 798
rect 1538 742 1550 798
rect 1470 708 1550 742
rect 1470 652 1482 708
rect 1538 652 1550 708
rect 1470 618 1550 652
rect 1470 562 1482 618
rect 1538 562 1550 618
rect 1470 528 1550 562
rect 1470 472 1482 528
rect 1538 472 1550 528
rect 1470 460 1550 472
rect 1870 798 1950 820
rect 1870 742 1882 798
rect 1938 742 1950 798
rect 1870 708 1950 742
rect 1870 652 1882 708
rect 1938 652 1950 708
rect 1870 618 1950 652
rect 1870 562 1882 618
rect 1938 562 1950 618
rect 1870 528 1950 562
rect 1870 472 1882 528
rect 1938 472 1950 528
rect 1870 460 1950 472
rect 2270 798 2350 820
rect 2270 742 2282 798
rect 2338 742 2350 798
rect 2270 708 2350 742
rect 2270 652 2282 708
rect 2338 652 2350 708
rect 2270 618 2350 652
rect 2270 562 2282 618
rect 2338 562 2350 618
rect 2270 528 2350 562
rect 2270 472 2282 528
rect 2338 472 2350 528
rect 2270 460 2350 472
rect 2670 798 2750 820
rect 2670 742 2682 798
rect 2738 742 2750 798
rect 2670 708 2750 742
rect 2670 652 2682 708
rect 2738 652 2750 708
rect 2670 618 2750 652
rect 2670 562 2682 618
rect 2738 562 2750 618
rect 2670 528 2750 562
rect 2670 472 2682 528
rect 2738 472 2750 528
rect 2670 460 2750 472
rect 3070 798 3150 820
rect 3070 742 3082 798
rect 3138 742 3150 798
rect 3070 708 3150 742
rect 3070 652 3082 708
rect 3138 652 3150 708
rect 3070 618 3150 652
rect 3070 562 3082 618
rect 3138 562 3150 618
rect 3070 528 3150 562
rect 3070 472 3082 528
rect 3138 472 3150 528
rect 3070 460 3150 472
rect 3470 798 3550 820
rect 3470 742 3482 798
rect 3538 742 3550 798
rect 3470 708 3550 742
rect 3470 652 3482 708
rect 3538 652 3550 708
rect 3470 618 3550 652
rect 3470 562 3482 618
rect 3538 562 3550 618
rect 3470 528 3550 562
rect 3470 472 3482 528
rect 3538 472 3550 528
rect 3470 460 3550 472
rect -60 176 20 180
rect -60 124 -46 176
rect 6 124 20 176
rect -60 100 20 124
rect -60 96 3840 100
rect -60 44 -46 96
rect 6 44 1294 96
rect 1346 44 1374 96
rect 1426 44 1694 96
rect 1746 44 1774 96
rect 1826 44 2094 96
rect 2146 44 2174 96
rect 2226 44 2494 96
rect 2546 44 2574 96
rect 2626 44 3840 96
rect -60 40 3840 44
rect 3980 86 4060 90
rect 3980 34 3994 86
rect 4046 34 4060 86
rect 3980 10 4060 34
rect 470 6 4060 10
rect 470 -46 494 6
rect 546 -46 574 6
rect 626 -46 894 6
rect 946 -46 974 6
rect 1026 -46 2894 6
rect 2946 -46 2974 6
rect 3026 -46 3294 6
rect 3346 -46 3374 6
rect 3426 -46 3994 6
rect 4046 -46 4060 6
rect 470 -50 4060 -46
<< via2 >>
rect -58 2942 -2 2998
rect 702 2792 758 2848
rect 792 2792 848 2848
rect 1052 2792 1108 2848
rect 1142 2792 1198 2848
rect 1452 2792 1508 2848
rect 1542 2792 1598 2848
rect 1852 2792 1908 2848
rect 1942 2792 1998 2848
rect 2252 2792 2308 2848
rect 2342 2792 2398 2848
rect 2652 2792 2708 2848
rect 2742 2792 2798 2848
rect 3052 2792 3108 2848
rect 3142 2792 3198 2848
rect 3452 2792 3508 2848
rect 3542 2792 3598 2848
rect 4182 2792 4238 2848
rect 682 2016 738 2018
rect 682 1964 684 2016
rect 684 1964 736 2016
rect 736 1964 738 2016
rect 682 1962 738 1964
rect 682 1926 738 1928
rect 682 1874 684 1926
rect 684 1874 736 1926
rect 736 1874 738 1926
rect 682 1872 738 1874
rect 682 1836 738 1838
rect 682 1784 684 1836
rect 684 1784 736 1836
rect 736 1784 738 1836
rect 682 1782 738 1784
rect 682 1746 738 1748
rect 682 1694 684 1746
rect 684 1694 736 1746
rect 736 1694 738 1746
rect 682 1692 738 1694
rect 1082 2016 1138 2018
rect 1082 1964 1084 2016
rect 1084 1964 1136 2016
rect 1136 1964 1138 2016
rect 1082 1962 1138 1964
rect 1082 1926 1138 1928
rect 1082 1874 1084 1926
rect 1084 1874 1136 1926
rect 1136 1874 1138 1926
rect 1082 1872 1138 1874
rect 1082 1836 1138 1838
rect 1082 1784 1084 1836
rect 1084 1784 1136 1836
rect 1136 1784 1138 1836
rect 1082 1782 1138 1784
rect 1082 1746 1138 1748
rect 1082 1694 1084 1746
rect 1084 1694 1136 1746
rect 1136 1694 1138 1746
rect 1082 1692 1138 1694
rect 1482 2016 1538 2018
rect 1482 1964 1484 2016
rect 1484 1964 1536 2016
rect 1536 1964 1538 2016
rect 1482 1962 1538 1964
rect 1482 1926 1538 1928
rect 1482 1874 1484 1926
rect 1484 1874 1536 1926
rect 1536 1874 1538 1926
rect 1482 1872 1538 1874
rect 1482 1836 1538 1838
rect 1482 1784 1484 1836
rect 1484 1784 1536 1836
rect 1536 1784 1538 1836
rect 1482 1782 1538 1784
rect 1482 1746 1538 1748
rect 1482 1694 1484 1746
rect 1484 1694 1536 1746
rect 1536 1694 1538 1746
rect 1482 1692 1538 1694
rect 1882 2016 1938 2018
rect 1882 1964 1884 2016
rect 1884 1964 1936 2016
rect 1936 1964 1938 2016
rect 1882 1962 1938 1964
rect 1882 1926 1938 1928
rect 1882 1874 1884 1926
rect 1884 1874 1936 1926
rect 1936 1874 1938 1926
rect 1882 1872 1938 1874
rect 1882 1836 1938 1838
rect 1882 1784 1884 1836
rect 1884 1784 1936 1836
rect 1936 1784 1938 1836
rect 1882 1782 1938 1784
rect 1882 1746 1938 1748
rect 1882 1694 1884 1746
rect 1884 1694 1936 1746
rect 1936 1694 1938 1746
rect 1882 1692 1938 1694
rect 2282 2016 2338 2018
rect 2282 1964 2284 2016
rect 2284 1964 2336 2016
rect 2336 1964 2338 2016
rect 2282 1962 2338 1964
rect 2282 1926 2338 1928
rect 2282 1874 2284 1926
rect 2284 1874 2336 1926
rect 2336 1874 2338 1926
rect 2282 1872 2338 1874
rect 2282 1836 2338 1838
rect 2282 1784 2284 1836
rect 2284 1784 2336 1836
rect 2336 1784 2338 1836
rect 2282 1782 2338 1784
rect 2282 1746 2338 1748
rect 2282 1694 2284 1746
rect 2284 1694 2336 1746
rect 2336 1694 2338 1746
rect 2282 1692 2338 1694
rect 2682 2016 2738 2018
rect 2682 1964 2684 2016
rect 2684 1964 2736 2016
rect 2736 1964 2738 2016
rect 2682 1962 2738 1964
rect 2682 1926 2738 1928
rect 2682 1874 2684 1926
rect 2684 1874 2736 1926
rect 2736 1874 2738 1926
rect 2682 1872 2738 1874
rect 2682 1836 2738 1838
rect 2682 1784 2684 1836
rect 2684 1784 2736 1836
rect 2736 1784 2738 1836
rect 2682 1782 2738 1784
rect 2682 1746 2738 1748
rect 2682 1694 2684 1746
rect 2684 1694 2736 1746
rect 2736 1694 2738 1746
rect 2682 1692 2738 1694
rect 3082 2016 3138 2018
rect 3082 1964 3084 2016
rect 3084 1964 3136 2016
rect 3136 1964 3138 2016
rect 3082 1962 3138 1964
rect 3082 1926 3138 1928
rect 3082 1874 3084 1926
rect 3084 1874 3136 1926
rect 3136 1874 3138 1926
rect 3082 1872 3138 1874
rect 3082 1836 3138 1838
rect 3082 1784 3084 1836
rect 3084 1784 3136 1836
rect 3136 1784 3138 1836
rect 3082 1782 3138 1784
rect 3082 1746 3138 1748
rect 3082 1694 3084 1746
rect 3084 1694 3136 1746
rect 3136 1694 3138 1746
rect 3082 1692 3138 1694
rect 3482 2016 3538 2018
rect 3482 1964 3484 2016
rect 3484 1964 3536 2016
rect 3536 1964 3538 2016
rect 3482 1962 3538 1964
rect 3482 1926 3538 1928
rect 3482 1874 3484 1926
rect 3484 1874 3536 1926
rect 3536 1874 3538 1926
rect 3482 1872 3538 1874
rect 3482 1836 3538 1838
rect 3482 1784 3484 1836
rect 3484 1784 3536 1836
rect 3536 1784 3538 1836
rect 3482 1782 3538 1784
rect 3482 1746 3538 1748
rect 3482 1694 3484 1746
rect 3484 1694 3536 1746
rect 3536 1694 3538 1746
rect 3482 1692 3538 1694
rect -168 1192 -112 1248
rect 682 796 738 798
rect 682 744 684 796
rect 684 744 736 796
rect 736 744 738 796
rect 682 742 738 744
rect 682 706 738 708
rect 682 654 684 706
rect 684 654 736 706
rect 736 654 738 706
rect 682 652 738 654
rect 682 616 738 618
rect 682 564 684 616
rect 684 564 736 616
rect 736 564 738 616
rect 682 562 738 564
rect 682 526 738 528
rect 682 474 684 526
rect 684 474 736 526
rect 736 474 738 526
rect 682 472 738 474
rect 1082 796 1138 798
rect 1082 744 1084 796
rect 1084 744 1136 796
rect 1136 744 1138 796
rect 1082 742 1138 744
rect 1082 706 1138 708
rect 1082 654 1084 706
rect 1084 654 1136 706
rect 1136 654 1138 706
rect 1082 652 1138 654
rect 1082 616 1138 618
rect 1082 564 1084 616
rect 1084 564 1136 616
rect 1136 564 1138 616
rect 1082 562 1138 564
rect 1082 526 1138 528
rect 1082 474 1084 526
rect 1084 474 1136 526
rect 1136 474 1138 526
rect 1082 472 1138 474
rect 1482 796 1538 798
rect 1482 744 1484 796
rect 1484 744 1536 796
rect 1536 744 1538 796
rect 1482 742 1538 744
rect 1482 706 1538 708
rect 1482 654 1484 706
rect 1484 654 1536 706
rect 1536 654 1538 706
rect 1482 652 1538 654
rect 1482 616 1538 618
rect 1482 564 1484 616
rect 1484 564 1536 616
rect 1536 564 1538 616
rect 1482 562 1538 564
rect 1482 526 1538 528
rect 1482 474 1484 526
rect 1484 474 1536 526
rect 1536 474 1538 526
rect 1482 472 1538 474
rect 1882 796 1938 798
rect 1882 744 1884 796
rect 1884 744 1936 796
rect 1936 744 1938 796
rect 1882 742 1938 744
rect 1882 706 1938 708
rect 1882 654 1884 706
rect 1884 654 1936 706
rect 1936 654 1938 706
rect 1882 652 1938 654
rect 1882 616 1938 618
rect 1882 564 1884 616
rect 1884 564 1936 616
rect 1936 564 1938 616
rect 1882 562 1938 564
rect 1882 526 1938 528
rect 1882 474 1884 526
rect 1884 474 1936 526
rect 1936 474 1938 526
rect 1882 472 1938 474
rect 2282 796 2338 798
rect 2282 744 2284 796
rect 2284 744 2336 796
rect 2336 744 2338 796
rect 2282 742 2338 744
rect 2282 706 2338 708
rect 2282 654 2284 706
rect 2284 654 2336 706
rect 2336 654 2338 706
rect 2282 652 2338 654
rect 2282 616 2338 618
rect 2282 564 2284 616
rect 2284 564 2336 616
rect 2336 564 2338 616
rect 2282 562 2338 564
rect 2282 526 2338 528
rect 2282 474 2284 526
rect 2284 474 2336 526
rect 2336 474 2338 526
rect 2282 472 2338 474
rect 2682 796 2738 798
rect 2682 744 2684 796
rect 2684 744 2736 796
rect 2736 744 2738 796
rect 2682 742 2738 744
rect 2682 706 2738 708
rect 2682 654 2684 706
rect 2684 654 2736 706
rect 2736 654 2738 706
rect 2682 652 2738 654
rect 2682 616 2738 618
rect 2682 564 2684 616
rect 2684 564 2736 616
rect 2736 564 2738 616
rect 2682 562 2738 564
rect 2682 526 2738 528
rect 2682 474 2684 526
rect 2684 474 2736 526
rect 2736 474 2738 526
rect 2682 472 2738 474
rect 3082 796 3138 798
rect 3082 744 3084 796
rect 3084 744 3136 796
rect 3136 744 3138 796
rect 3082 742 3138 744
rect 3082 706 3138 708
rect 3082 654 3084 706
rect 3084 654 3136 706
rect 3136 654 3138 706
rect 3082 652 3138 654
rect 3082 616 3138 618
rect 3082 564 3084 616
rect 3084 564 3136 616
rect 3136 564 3138 616
rect 3082 562 3138 564
rect 3082 526 3138 528
rect 3082 474 3084 526
rect 3084 474 3136 526
rect 3136 474 3138 526
rect 3082 472 3138 474
rect 3482 796 3538 798
rect 3482 744 3484 796
rect 3484 744 3536 796
rect 3536 744 3538 796
rect 3482 742 3538 744
rect 3482 706 3538 708
rect 3482 654 3484 706
rect 3484 654 3536 706
rect 3536 654 3538 706
rect 3482 652 3538 654
rect 3482 616 3538 618
rect 3482 564 3484 616
rect 3484 564 3536 616
rect 3536 564 3538 616
rect 3482 562 3538 564
rect 3482 526 3538 528
rect 3482 474 3484 526
rect 3484 474 3536 526
rect 3536 474 3538 526
rect 3482 472 3538 474
<< metal3 >>
rect -280 2920 -180 3020
rect -80 2998 20 3020
rect -80 2942 -58 2998
rect -2 2942 20 2998
rect -80 2920 20 2942
rect -270 2860 -190 2920
rect -270 2780 -100 2860
rect -180 1248 -100 2780
rect 690 2848 860 2860
rect 690 2792 702 2848
rect 758 2792 792 2848
rect 848 2792 860 2848
rect 690 2780 860 2792
rect 1040 2848 1210 2860
rect 1040 2792 1052 2848
rect 1108 2792 1142 2848
rect 1198 2792 1210 2848
rect 1040 2780 1210 2792
rect 1440 2848 1610 2860
rect 1440 2792 1452 2848
rect 1508 2792 1542 2848
rect 1598 2792 1610 2848
rect 1440 2780 1610 2792
rect 1840 2848 2010 2860
rect 1840 2792 1852 2848
rect 1908 2792 1942 2848
rect 1998 2792 2010 2848
rect 1840 2780 2010 2792
rect 2240 2848 2410 2860
rect 2240 2792 2252 2848
rect 2308 2792 2342 2848
rect 2398 2792 2410 2848
rect 2240 2780 2410 2792
rect 2640 2848 2810 2860
rect 2640 2792 2652 2848
rect 2708 2792 2742 2848
rect 2798 2792 2810 2848
rect 2640 2780 2810 2792
rect 3040 2848 3210 2860
rect 3040 2792 3052 2848
rect 3108 2792 3142 2848
rect 3198 2792 3210 2848
rect 3040 2780 3210 2792
rect 3440 2848 3610 2860
rect 3440 2792 3452 2848
rect 3508 2792 3542 2848
rect 3598 2792 3610 2848
rect 3440 2780 3610 2792
rect 4160 2848 4260 2870
rect 4160 2792 4182 2848
rect 4238 2792 4260 2848
rect 690 2040 750 2780
rect 1090 2040 1150 2780
rect 1490 2040 1550 2780
rect 1890 2040 1950 2780
rect 2290 2040 2350 2780
rect 2690 2040 2750 2780
rect 3090 2040 3150 2780
rect 3490 2040 3550 2780
rect 4160 2770 4260 2792
rect 670 2018 750 2040
rect 670 1962 682 2018
rect 738 1962 750 2018
rect 670 1928 750 1962
rect 670 1872 682 1928
rect 738 1872 750 1928
rect 670 1838 750 1872
rect 670 1782 682 1838
rect 738 1782 750 1838
rect 670 1748 750 1782
rect 670 1692 682 1748
rect 738 1692 750 1748
rect 670 1680 750 1692
rect 1070 2018 1150 2040
rect 1070 1962 1082 2018
rect 1138 1962 1150 2018
rect 1070 1928 1150 1962
rect 1070 1872 1082 1928
rect 1138 1872 1150 1928
rect 1070 1838 1150 1872
rect 1070 1782 1082 1838
rect 1138 1782 1150 1838
rect 1070 1748 1150 1782
rect 1070 1692 1082 1748
rect 1138 1692 1150 1748
rect 1070 1680 1150 1692
rect 1470 2018 1550 2040
rect 1470 1962 1482 2018
rect 1538 1962 1550 2018
rect 1470 1928 1550 1962
rect 1470 1872 1482 1928
rect 1538 1872 1550 1928
rect 1470 1838 1550 1872
rect 1470 1782 1482 1838
rect 1538 1782 1550 1838
rect 1470 1748 1550 1782
rect 1470 1692 1482 1748
rect 1538 1692 1550 1748
rect 1470 1680 1550 1692
rect 1870 2018 1950 2040
rect 1870 1962 1882 2018
rect 1938 1962 1950 2018
rect 1870 1928 1950 1962
rect 1870 1872 1882 1928
rect 1938 1872 1950 1928
rect 1870 1838 1950 1872
rect 1870 1782 1882 1838
rect 1938 1782 1950 1838
rect 1870 1748 1950 1782
rect 1870 1692 1882 1748
rect 1938 1692 1950 1748
rect 1870 1680 1950 1692
rect 2270 2018 2350 2040
rect 2270 1962 2282 2018
rect 2338 1962 2350 2018
rect 2270 1928 2350 1962
rect 2270 1872 2282 1928
rect 2338 1872 2350 1928
rect 2270 1838 2350 1872
rect 2270 1782 2282 1838
rect 2338 1782 2350 1838
rect 2270 1748 2350 1782
rect 2270 1692 2282 1748
rect 2338 1692 2350 1748
rect 2270 1680 2350 1692
rect 2670 2018 2750 2040
rect 2670 1962 2682 2018
rect 2738 1962 2750 2018
rect 2670 1928 2750 1962
rect 2670 1872 2682 1928
rect 2738 1872 2750 1928
rect 2670 1838 2750 1872
rect 2670 1782 2682 1838
rect 2738 1782 2750 1838
rect 2670 1748 2750 1782
rect 2670 1692 2682 1748
rect 2738 1692 2750 1748
rect 2670 1680 2750 1692
rect 3070 2018 3150 2040
rect 3070 1962 3082 2018
rect 3138 1962 3150 2018
rect 3070 1928 3150 1962
rect 3070 1872 3082 1928
rect 3138 1872 3150 1928
rect 3070 1838 3150 1872
rect 3070 1782 3082 1838
rect 3138 1782 3150 1838
rect 3070 1748 3150 1782
rect 3070 1692 3082 1748
rect 3138 1692 3150 1748
rect 3070 1680 3150 1692
rect 3470 2018 3550 2040
rect 3470 1962 3482 2018
rect 3538 1962 3550 2018
rect 3470 1928 3550 1962
rect 3470 1872 3482 1928
rect 3538 1872 3550 1928
rect 3470 1838 3550 1872
rect 3470 1782 3482 1838
rect 3538 1782 3550 1838
rect 3470 1748 3550 1782
rect 3470 1692 3482 1748
rect 3538 1692 3550 1748
rect 3470 1680 3550 1692
rect -180 1192 -168 1248
rect -112 1192 -100 1248
rect -180 1180 -100 1192
rect 690 820 750 1680
rect 1090 820 1150 1680
rect 1490 820 1550 1680
rect 1890 820 1950 1680
rect 2290 820 2350 1680
rect 2690 820 2750 1680
rect 3090 820 3150 1680
rect 3490 820 3550 1680
rect 670 798 750 820
rect 670 742 682 798
rect 738 742 750 798
rect 670 708 750 742
rect 670 652 682 708
rect 738 652 750 708
rect 670 618 750 652
rect 670 562 682 618
rect 738 562 750 618
rect 670 528 750 562
rect 670 472 682 528
rect 738 472 750 528
rect 670 460 750 472
rect 1070 798 1150 820
rect 1070 742 1082 798
rect 1138 742 1150 798
rect 1070 708 1150 742
rect 1070 652 1082 708
rect 1138 652 1150 708
rect 1070 618 1150 652
rect 1070 562 1082 618
rect 1138 562 1150 618
rect 1070 528 1150 562
rect 1070 472 1082 528
rect 1138 472 1150 528
rect 1070 460 1150 472
rect 1470 798 1550 820
rect 1470 742 1482 798
rect 1538 742 1550 798
rect 1470 708 1550 742
rect 1470 652 1482 708
rect 1538 652 1550 708
rect 1470 618 1550 652
rect 1470 562 1482 618
rect 1538 562 1550 618
rect 1470 528 1550 562
rect 1470 472 1482 528
rect 1538 472 1550 528
rect 1470 460 1550 472
rect 1870 798 1950 820
rect 1870 742 1882 798
rect 1938 742 1950 798
rect 1870 708 1950 742
rect 1870 652 1882 708
rect 1938 652 1950 708
rect 1870 618 1950 652
rect 1870 562 1882 618
rect 1938 562 1950 618
rect 1870 528 1950 562
rect 1870 472 1882 528
rect 1938 472 1950 528
rect 1870 460 1950 472
rect 2270 798 2350 820
rect 2270 742 2282 798
rect 2338 742 2350 798
rect 2270 708 2350 742
rect 2270 652 2282 708
rect 2338 652 2350 708
rect 2270 618 2350 652
rect 2270 562 2282 618
rect 2338 562 2350 618
rect 2270 528 2350 562
rect 2270 472 2282 528
rect 2338 472 2350 528
rect 2270 460 2350 472
rect 2670 798 2750 820
rect 2670 742 2682 798
rect 2738 742 2750 798
rect 2670 708 2750 742
rect 2670 652 2682 708
rect 2738 652 2750 708
rect 2670 618 2750 652
rect 2670 562 2682 618
rect 2738 562 2750 618
rect 2670 528 2750 562
rect 2670 472 2682 528
rect 2738 472 2750 528
rect 2670 460 2750 472
rect 3070 798 3150 820
rect 3070 742 3082 798
rect 3138 742 3150 798
rect 3070 708 3150 742
rect 3070 652 3082 708
rect 3138 652 3150 708
rect 3070 618 3150 652
rect 3070 562 3082 618
rect 3138 562 3150 618
rect 3070 528 3150 562
rect 3070 472 3082 528
rect 3138 472 3150 528
rect 3070 460 3150 472
rect 3470 798 3550 820
rect 3470 742 3482 798
rect 3538 742 3550 798
rect 3470 708 3550 742
rect 3470 652 3482 708
rect 3538 652 3550 708
rect 3470 618 3550 652
rect 3470 562 3482 618
rect 3538 562 3550 618
rect 3470 528 3550 562
rect 3470 472 3482 528
rect 3538 472 3550 528
rect 3470 460 3550 472
rect 690 240 750 460
rect 1090 240 1150 460
rect 1490 240 1550 460
rect 1890 240 1950 460
rect 2290 240 2350 460
rect 2690 240 2750 460
rect 3090 240 3150 460
rect 3490 240 3550 460
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_0
timestamp 1757161594
transform 0 1 3798 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_1
timestamp 1757161594
transform 0 1 2598 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_2
timestamp 1757161594
transform 0 1 2998 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_3
timestamp 1757161594
transform 0 1 998 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_4
timestamp 1757161594
transform 0 1 598 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_5
timestamp 1757161594
transform 0 1 198 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_6
timestamp 1757161594
transform 0 1 1398 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_7
timestamp 1757161594
transform 0 1 1798 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_8
timestamp 1757161594
transform 0 1 2198 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_9
timestamp 1757161594
transform 0 1 3398 1 0 594
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_10
timestamp 1757161594
transform 0 1 3798 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_11
timestamp 1757161594
transform 0 1 3398 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_12
timestamp 1757161594
transform 0 1 2998 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_13
timestamp 1757161594
transform 0 1 2598 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_14
timestamp 1757161594
transform 0 1 2198 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_15
timestamp 1757161594
transform 0 1 1798 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_16
timestamp 1757161594
transform 0 1 1398 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_17
timestamp 1757161594
transform 0 1 998 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_18
timestamp 1757161594
transform 0 1 598 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_21
timestamp 1757161594
transform 0 1 198 1 0 1824
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_0
timestamp 1757161594
transform 0 1 1398 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_1
timestamp 1757161594
transform 0 1 598 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_2
timestamp 1757161594
transform 0 1 998 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_3
timestamp 1757161594
transform 0 1 198 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_4
timestamp 1757161594
transform 0 1 1798 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_5
timestamp 1757161594
transform 0 1 2198 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_6
timestamp 1757161594
transform 0 1 2598 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_7
timestamp 1757161594
transform 0 1 2998 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_8
timestamp 1757161594
transform 0 1 3398 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_9
timestamp 1757161594
transform 0 1 3798 1 0 -236
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_12
timestamp 1757161594
transform 0 1 198 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_13
timestamp 1757161594
transform 0 1 1398 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_14
timestamp 1757161594
transform 0 1 2198 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_15
timestamp 1757161594
transform 0 1 1798 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_16
timestamp 1757161594
transform 0 1 2998 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_17
timestamp 1757161594
transform 0 1 2598 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_18
timestamp 1757161594
transform 0 1 3398 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_19
timestamp 1757161594
transform 0 1 598 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_20
timestamp 1757161594
transform 0 1 3798 1 0 2614
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_21
timestamp 1757161594
transform 0 1 998 1 0 2614
box -194 -198 194 164
<< labels >>
flabel metal3 s 4160 2770 4260 2870 0 FreeSans 782 0 0 0 Vin
port 0 nsew
<< end >>
