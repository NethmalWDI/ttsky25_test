magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< error_s >>
rect 368 -437 556 -424
rect 400 -473 654 -460
rect 520 -500 654 -473
rect 1690 -560 1778 -500
<< nwell >>
rect -80 -460 2530 2710
rect -80 -500 400 -460
rect 520 -500 2530 -460
rect 1610 -560 1690 -500
<< nsubdiff >>
rect 3 2593 96 2627
rect 130 2593 164 2627
rect 198 2593 232 2627
rect 266 2593 300 2627
rect 334 2593 368 2627
rect 402 2593 436 2627
rect 470 2593 504 2627
rect 538 2593 572 2627
rect 606 2593 640 2627
rect 674 2593 708 2627
rect 742 2593 776 2627
rect 810 2593 844 2627
rect 878 2593 912 2627
rect 946 2593 980 2627
rect 1014 2593 1048 2627
rect 1082 2593 1116 2627
rect 1150 2593 1184 2627
rect 1218 2593 1252 2627
rect 1286 2593 1320 2627
rect 1354 2593 1388 2627
rect 1422 2593 1456 2627
rect 1490 2593 1524 2627
rect 1558 2593 1592 2627
rect 1626 2593 1660 2627
rect 1694 2593 1728 2627
rect 1762 2593 1796 2627
rect 1830 2593 1864 2627
rect 1898 2593 1932 2627
rect 1966 2593 2000 2627
rect 2034 2593 2068 2627
rect 2102 2593 2136 2627
rect 2170 2593 2204 2627
rect 2238 2593 2272 2627
rect 2306 2593 2340 2627
rect 2374 2593 2467 2627
rect 3 2545 37 2593
rect 3 2477 37 2511
rect 3 2409 37 2443
rect 3 2341 37 2375
rect 3 2273 37 2307
rect 3 2205 37 2239
rect 3 2137 37 2171
rect 3 2069 37 2103
rect 3 2001 37 2035
rect 3 1933 37 1967
rect 3 1865 37 1899
rect 3 1797 37 1831
rect 3 1729 37 1763
rect 3 1661 37 1695
rect 3 1593 37 1627
rect 3 1525 37 1559
rect 3 1457 37 1491
rect 3 1389 37 1423
rect 3 1321 37 1355
rect 3 1253 37 1287
rect 3 1185 37 1219
rect 3 1117 37 1151
rect 3 1049 37 1083
rect 3 981 37 1015
rect 3 913 37 947
rect 3 845 37 879
rect 3 777 37 811
rect 3 709 37 743
rect 3 641 37 675
rect 3 573 37 607
rect 3 505 37 539
rect 3 437 37 471
rect 3 369 37 403
rect 3 301 37 335
rect 3 233 37 267
rect 3 165 37 199
rect 3 97 37 131
rect 3 29 37 63
rect 3 -39 37 -5
rect 3 -107 37 -73
rect 3 -175 37 -141
rect 3 -243 37 -209
rect 3 -311 37 -277
rect 3 -403 37 -345
rect 2433 2545 2467 2593
rect 2433 2477 2467 2511
rect 2433 2409 2467 2443
rect 2433 2341 2467 2375
rect 2433 2273 2467 2307
rect 2433 2205 2467 2239
rect 2433 2137 2467 2171
rect 2433 2069 2467 2103
rect 2433 2001 2467 2035
rect 2433 1933 2467 1967
rect 2433 1865 2467 1899
rect 2433 1797 2467 1831
rect 2433 1729 2467 1763
rect 2433 1661 2467 1695
rect 2433 1593 2467 1627
rect 2433 1525 2467 1559
rect 2433 1457 2467 1491
rect 2433 1389 2467 1423
rect 2433 1321 2467 1355
rect 2433 1253 2467 1287
rect 2433 1185 2467 1219
rect 2433 1117 2467 1151
rect 2433 1049 2467 1083
rect 2433 981 2467 1015
rect 2433 913 2467 947
rect 2433 845 2467 879
rect 2433 777 2467 811
rect 2433 709 2467 743
rect 2433 641 2467 675
rect 2433 573 2467 607
rect 2433 505 2467 539
rect 2433 437 2467 471
rect 2433 369 2467 403
rect 2433 301 2467 335
rect 2433 233 2467 267
rect 2433 165 2467 199
rect 2433 97 2467 131
rect 2433 29 2467 63
rect 2433 -39 2467 -5
rect 2433 -107 2467 -73
rect 2433 -175 2467 -141
rect 2433 -243 2467 -209
rect 2433 -311 2467 -277
rect 2433 -403 2467 -345
rect 3 -437 96 -403
rect 130 -437 164 -403
rect 198 -437 232 -403
rect 266 -437 300 -403
rect 334 -437 368 -403
rect 402 -437 436 -403
rect 470 -437 504 -403
rect 538 -437 572 -403
rect 606 -437 640 -403
rect 674 -437 708 -403
rect 742 -437 776 -403
rect 810 -437 844 -403
rect 878 -437 912 -403
rect 946 -437 980 -403
rect 1014 -437 1048 -403
rect 1082 -437 1116 -403
rect 1150 -437 1184 -403
rect 1218 -437 1252 -403
rect 1286 -437 1320 -403
rect 1354 -437 1388 -403
rect 1422 -437 1456 -403
rect 1490 -437 1524 -403
rect 1558 -437 1592 -403
rect 1626 -437 1660 -403
rect 1694 -437 1728 -403
rect 1762 -437 1796 -403
rect 1830 -437 1864 -403
rect 1898 -437 1932 -403
rect 1966 -437 2000 -403
rect 2034 -437 2068 -403
rect 2102 -437 2136 -403
rect 2170 -437 2204 -403
rect 2238 -437 2272 -403
rect 2306 -437 2340 -403
rect 2374 -437 2467 -403
<< nsubdiffcont >>
rect 96 2593 130 2627
rect 164 2593 198 2627
rect 232 2593 266 2627
rect 300 2593 334 2627
rect 368 2593 402 2627
rect 436 2593 470 2627
rect 504 2593 538 2627
rect 572 2593 606 2627
rect 640 2593 674 2627
rect 708 2593 742 2627
rect 776 2593 810 2627
rect 844 2593 878 2627
rect 912 2593 946 2627
rect 980 2593 1014 2627
rect 1048 2593 1082 2627
rect 1116 2593 1150 2627
rect 1184 2593 1218 2627
rect 1252 2593 1286 2627
rect 1320 2593 1354 2627
rect 1388 2593 1422 2627
rect 1456 2593 1490 2627
rect 1524 2593 1558 2627
rect 1592 2593 1626 2627
rect 1660 2593 1694 2627
rect 1728 2593 1762 2627
rect 1796 2593 1830 2627
rect 1864 2593 1898 2627
rect 1932 2593 1966 2627
rect 2000 2593 2034 2627
rect 2068 2593 2102 2627
rect 2136 2593 2170 2627
rect 2204 2593 2238 2627
rect 2272 2593 2306 2627
rect 2340 2593 2374 2627
rect 3 2511 37 2545
rect 3 2443 37 2477
rect 3 2375 37 2409
rect 3 2307 37 2341
rect 3 2239 37 2273
rect 3 2171 37 2205
rect 3 2103 37 2137
rect 3 2035 37 2069
rect 3 1967 37 2001
rect 3 1899 37 1933
rect 3 1831 37 1865
rect 3 1763 37 1797
rect 3 1695 37 1729
rect 3 1627 37 1661
rect 3 1559 37 1593
rect 3 1491 37 1525
rect 3 1423 37 1457
rect 3 1355 37 1389
rect 3 1287 37 1321
rect 3 1219 37 1253
rect 3 1151 37 1185
rect 3 1083 37 1117
rect 3 1015 37 1049
rect 3 947 37 981
rect 3 879 37 913
rect 3 811 37 845
rect 3 743 37 777
rect 3 675 37 709
rect 3 607 37 641
rect 3 539 37 573
rect 3 471 37 505
rect 3 403 37 437
rect 3 335 37 369
rect 3 267 37 301
rect 3 199 37 233
rect 3 131 37 165
rect 3 63 37 97
rect 3 -5 37 29
rect 3 -73 37 -39
rect 3 -141 37 -107
rect 3 -209 37 -175
rect 3 -277 37 -243
rect 3 -345 37 -311
rect 2433 2511 2467 2545
rect 2433 2443 2467 2477
rect 2433 2375 2467 2409
rect 2433 2307 2467 2341
rect 2433 2239 2467 2273
rect 2433 2171 2467 2205
rect 2433 2103 2467 2137
rect 2433 2035 2467 2069
rect 2433 1967 2467 2001
rect 2433 1899 2467 1933
rect 2433 1831 2467 1865
rect 2433 1763 2467 1797
rect 2433 1695 2467 1729
rect 2433 1627 2467 1661
rect 2433 1559 2467 1593
rect 2433 1491 2467 1525
rect 2433 1423 2467 1457
rect 2433 1355 2467 1389
rect 2433 1287 2467 1321
rect 2433 1219 2467 1253
rect 2433 1151 2467 1185
rect 2433 1083 2467 1117
rect 2433 1015 2467 1049
rect 2433 947 2467 981
rect 2433 879 2467 913
rect 2433 811 2467 845
rect 2433 743 2467 777
rect 2433 675 2467 709
rect 2433 607 2467 641
rect 2433 539 2467 573
rect 2433 471 2467 505
rect 2433 403 2467 437
rect 2433 335 2467 369
rect 2433 267 2467 301
rect 2433 199 2467 233
rect 2433 131 2467 165
rect 2433 63 2467 97
rect 2433 -5 2467 29
rect 2433 -73 2467 -39
rect 2433 -141 2467 -107
rect 2433 -209 2467 -175
rect 2433 -277 2467 -243
rect 2433 -345 2467 -311
rect 96 -437 130 -403
rect 164 -437 198 -403
rect 232 -437 266 -403
rect 300 -437 334 -403
rect 368 -437 402 -403
rect 436 -437 470 -403
rect 504 -437 538 -403
rect 572 -437 606 -403
rect 640 -437 674 -403
rect 708 -437 742 -403
rect 776 -437 810 -403
rect 844 -437 878 -403
rect 912 -437 946 -403
rect 980 -437 1014 -403
rect 1048 -437 1082 -403
rect 1116 -437 1150 -403
rect 1184 -437 1218 -403
rect 1252 -437 1286 -403
rect 1320 -437 1354 -403
rect 1388 -437 1422 -403
rect 1456 -437 1490 -403
rect 1524 -437 1558 -403
rect 1592 -437 1626 -403
rect 1660 -437 1694 -403
rect 1728 -437 1762 -403
rect 1796 -437 1830 -403
rect 1864 -437 1898 -403
rect 1932 -437 1966 -403
rect 2000 -437 2034 -403
rect 2068 -437 2102 -403
rect 2136 -437 2170 -403
rect 2204 -437 2238 -403
rect 2272 -437 2306 -403
rect 2340 -437 2374 -403
<< locali >>
rect 3 2593 96 2627
rect 130 2593 164 2627
rect 198 2593 232 2627
rect 266 2593 300 2627
rect 334 2593 368 2627
rect 402 2593 436 2627
rect 470 2593 504 2627
rect 538 2593 572 2627
rect 606 2593 640 2627
rect 674 2593 708 2627
rect 742 2593 776 2627
rect 810 2593 844 2627
rect 878 2593 912 2627
rect 946 2593 980 2627
rect 1014 2593 1048 2627
rect 1082 2593 1116 2627
rect 1150 2593 1184 2627
rect 1218 2593 1252 2627
rect 1286 2593 1320 2627
rect 1354 2593 1388 2627
rect 1422 2593 1456 2627
rect 1490 2593 1524 2627
rect 1558 2593 1592 2627
rect 1626 2593 1660 2627
rect 1694 2593 1728 2627
rect 1762 2593 1796 2627
rect 1830 2593 1864 2627
rect 1898 2593 1932 2627
rect 1966 2593 2000 2627
rect 2034 2593 2068 2627
rect 2102 2593 2136 2627
rect 2170 2593 2204 2627
rect 2238 2593 2272 2627
rect 2306 2593 2340 2627
rect 2374 2593 2467 2627
rect 3 2545 37 2593
rect 3 2477 37 2511
rect 3 2409 37 2443
rect 3 2341 37 2375
rect 3 2273 37 2307
rect 3 2205 37 2239
rect 3 2137 37 2171
rect 3 2069 37 2103
rect 3 2001 37 2035
rect 3 1933 37 1967
rect 3 1865 37 1899
rect 3 1797 37 1831
rect 3 1729 37 1763
rect 3 1661 37 1695
rect 3 1593 37 1627
rect 3 1525 37 1559
rect 3 1457 37 1491
rect 3 1389 37 1423
rect 3 1321 37 1355
rect 3 1253 37 1287
rect 3 1185 37 1219
rect 3 1117 37 1151
rect 3 1049 37 1083
rect 3 981 37 1015
rect 3 913 37 947
rect 3 845 37 879
rect 3 777 37 811
rect 3 709 37 743
rect 3 641 37 675
rect 3 573 37 607
rect 3 505 37 539
rect 3 437 37 471
rect 3 369 37 403
rect 3 301 37 335
rect 3 233 37 267
rect 3 165 37 199
rect 3 97 37 131
rect 3 29 37 63
rect 3 -39 37 -5
rect 3 -107 37 -73
rect 3 -175 37 -141
rect 3 -243 37 -209
rect 3 -311 37 -277
rect 3 -403 37 -345
rect 2433 2545 2467 2593
rect 2433 2477 2467 2511
rect 2433 2409 2467 2443
rect 2433 2341 2467 2375
rect 2433 2273 2467 2307
rect 2433 2205 2467 2239
rect 2433 2137 2467 2171
rect 2433 2069 2467 2103
rect 2433 2001 2467 2035
rect 2433 1933 2467 1967
rect 2433 1865 2467 1899
rect 2433 1797 2467 1831
rect 2433 1729 2467 1763
rect 2433 1661 2467 1695
rect 2433 1593 2467 1627
rect 2433 1525 2467 1559
rect 2433 1457 2467 1491
rect 2433 1389 2467 1423
rect 2433 1321 2467 1355
rect 2433 1253 2467 1287
rect 2433 1185 2467 1219
rect 2433 1117 2467 1151
rect 2433 1049 2467 1083
rect 2433 981 2467 1015
rect 2433 913 2467 947
rect 2433 845 2467 879
rect 2433 777 2467 811
rect 2433 709 2467 743
rect 2433 641 2467 675
rect 2433 573 2467 607
rect 2433 505 2467 539
rect 2433 437 2467 471
rect 2433 369 2467 403
rect 2433 301 2467 335
rect 2433 233 2467 267
rect 2433 165 2467 199
rect 2433 97 2467 131
rect 2433 29 2467 63
rect 2433 -39 2467 -5
rect 2433 -107 2467 -73
rect 2433 -175 2467 -141
rect 2433 -243 2467 -209
rect 2433 -311 2467 -277
rect 2433 -403 2467 -345
rect 3 -437 96 -403
rect 130 -437 164 -403
rect 198 -437 232 -403
rect 266 -437 300 -403
rect 334 -437 368 -403
rect 402 -437 436 -403
rect 470 -437 504 -403
rect 538 -437 572 -403
rect 606 -437 640 -403
rect 674 -437 708 -403
rect 742 -437 776 -403
rect 810 -437 844 -403
rect 878 -437 912 -403
rect 946 -437 980 -403
rect 1014 -437 1048 -403
rect 1082 -437 1116 -403
rect 1150 -437 1184 -403
rect 1218 -437 1252 -403
rect 1286 -437 1320 -403
rect 1354 -437 1388 -403
rect 1422 -437 1456 -403
rect 1490 -437 1524 -403
rect 1558 -437 1592 -403
rect 1626 -437 1660 -403
rect 1694 -437 1728 -403
rect 1762 -437 1796 -403
rect 1830 -437 1864 -403
rect 1898 -437 1932 -403
rect 1966 -437 2000 -403
rect 2034 -437 2068 -403
rect 2102 -437 2136 -403
rect 2170 -437 2204 -403
rect 2238 -437 2272 -403
rect 2306 -437 2340 -403
rect 2374 -437 2467 -403
<< metal1 >>
rect 110 2090 2390 2530
rect 330 90 390 2090
rect 100 -30 390 90
rect 480 96 680 100
rect 480 44 534 96
rect 586 44 614 96
rect 666 44 680 96
rect 480 40 680 44
rect 730 90 790 1800
rect 1130 90 1190 1800
rect 1530 240 1590 1800
rect 1930 240 1990 1800
rect 1510 226 1590 240
rect 1510 174 1524 226
rect 1576 174 1590 226
rect 1510 160 1590 174
rect 1910 226 1990 240
rect 1910 174 1924 226
rect 1976 174 1990 226
rect 1910 160 1990 174
rect 1530 90 1590 160
rect 730 40 1590 90
rect 1720 96 1880 100
rect 1720 44 1734 96
rect 1786 44 1814 96
rect 1866 44 1880 96
rect 1930 90 1990 160
rect 2330 90 2390 2090
rect 1720 40 1880 44
rect 2120 -30 2390 90
rect 100 -80 2390 -30
rect 110 -90 2390 -80
rect 120 -340 2390 -90
<< via1 >>
rect 534 44 586 96
rect 614 44 666 96
rect 1524 174 1576 226
rect 1924 174 1976 226
rect 1734 44 1786 96
rect 1814 44 1866 96
<< metal2 >>
rect 1510 228 1590 240
rect 1510 172 1522 228
rect 1578 172 1590 228
rect 1510 160 1590 172
rect 1910 228 1990 240
rect 1910 172 1922 228
rect 1978 172 1990 228
rect 1910 160 1990 172
rect 420 96 1880 100
rect 420 44 534 96
rect 586 44 614 96
rect 666 44 1734 96
rect 1786 44 1814 96
rect 1866 44 1880 96
rect 420 40 1880 44
rect 420 -450 480 40
rect 1610 -332 1690 -320
rect 1610 -388 1622 -332
rect 1678 -340 1690 -332
rect 1990 -332 2070 -320
rect 1990 -340 2002 -332
rect 1678 -388 2002 -340
rect 2058 -388 2070 -332
rect 1610 -410 2070 -388
rect 400 -482 520 -450
rect 400 -538 432 -482
rect 488 -538 520 -482
rect 400 -570 520 -538
<< via2 >>
rect 1522 226 1578 228
rect 1522 174 1524 226
rect 1524 174 1576 226
rect 1576 174 1578 226
rect 1522 172 1578 174
rect 1922 226 1978 228
rect 1922 174 1924 226
rect 1924 174 1976 226
rect 1976 174 1978 226
rect 1922 172 1978 174
rect 1622 -388 1678 -332
rect 2002 -388 2058 -332
rect 432 -538 488 -482
<< metal3 >>
rect 1510 228 1670 240
rect 1510 172 1522 228
rect 1578 172 1670 228
rect 1510 160 1670 172
rect 1910 228 2070 240
rect 1910 172 1922 228
rect 1978 172 2070 228
rect 1910 160 2070 172
rect 1610 -320 1670 160
rect 2010 -320 2070 160
rect 1610 -332 1690 -320
rect 1610 -388 1622 -332
rect 1678 -388 1690 -332
rect 400 -482 520 -450
rect 400 -538 432 -482
rect 488 -538 520 -482
rect 400 -570 520 -538
rect 1610 -560 1690 -388
rect 1990 -332 2070 -320
rect 1990 -388 2002 -332
rect 2058 -388 2070 -332
rect 1990 -410 2070 -388
use sky130_fd_pr__pfet_01v8_lvt_76U4T2  sky130_fd_pr__pfet_01v8_lvt_76U4T2_0
timestamp 1757161594
transform 0 1 2238 -1 0 1094
box -1094 -198 1094 164
use sky130_fd_pr__pfet_01v8_lvt_76U4T2  sky130_fd_pr__pfet_01v8_lvt_76U4T2_1
timestamp 1757161594
transform 0 1 1838 -1 0 1094
box -1094 -198 1094 164
use sky130_fd_pr__pfet_01v8_lvt_76U4T2  sky130_fd_pr__pfet_01v8_lvt_76U4T2_2
timestamp 1757161594
transform 0 1 638 -1 0 1094
box -1094 -198 1094 164
use sky130_fd_pr__pfet_01v8_lvt_76U4T2  sky130_fd_pr__pfet_01v8_lvt_76U4T2_4
timestamp 1757161594
transform 0 1 1038 -1 0 1094
box -1094 -198 1094 164
use sky130_fd_pr__pfet_01v8_lvt_76U4T2  sky130_fd_pr__pfet_01v8_lvt_76U4T2_5
timestamp 1757161594
transform 0 1 1438 -1 0 1094
box -1094 -198 1094 164
use sky130_fd_pr__pfet_01v8_lvt_76U4T2  sky130_fd_pr__pfet_01v8_lvt_76U4T2_6
timestamp 1757161594
transform 0 1 238 -1 0 1094
box -1094 -198 1094 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_0
timestamp 1757161594
transform 0 1 1438 -1 0 -186
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_1
timestamp 1757161594
transform 0 1 1038 -1 0 -186
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_2
timestamp 1757161594
transform 0 1 638 -1 0 -186
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_3
timestamp 1757161594
transform 0 1 238 -1 0 -186
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_4
timestamp 1757161594
transform 0 1 1838 -1 0 -186
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_5
timestamp 1757161594
transform 0 1 2238 -1 0 -186
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_6
timestamp 1757161594
transform 0 1 238 -1 0 2374
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_7
timestamp 1757161594
transform 0 1 638 -1 0 2374
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_8
timestamp 1757161594
transform 0 1 1038 -1 0 2374
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_9
timestamp 1757161594
transform 0 1 1438 -1 0 2374
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_10
timestamp 1757161594
transform 0 1 1838 -1 0 2374
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_KVZWZ9  sky130_fd_pr__pfet_01v8_lvt_KVZWZ9_11
timestamp 1757161594
transform 0 1 2238 -1 0 2374
box -194 -198 194 164
<< end >>
