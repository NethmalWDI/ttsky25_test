magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< metal3 >>
rect -686 512 686 540
rect -686 448 602 512
rect 666 448 686 512
rect -686 432 686 448
rect -686 368 602 432
rect 666 368 686 432
rect -686 352 686 368
rect -686 288 602 352
rect 666 288 686 352
rect -686 272 686 288
rect -686 208 602 272
rect 666 208 686 272
rect -686 192 686 208
rect -686 128 602 192
rect 666 128 686 192
rect -686 112 686 128
rect -686 48 602 112
rect 666 48 686 112
rect -686 32 686 48
rect -686 -32 602 32
rect 666 -32 686 32
rect -686 -48 686 -32
rect -686 -112 602 -48
rect 666 -112 686 -48
rect -686 -128 686 -112
rect -686 -192 602 -128
rect 666 -192 686 -128
rect -686 -208 686 -192
rect -686 -272 602 -208
rect 666 -272 686 -208
rect -686 -288 686 -272
rect -686 -352 602 -288
rect 666 -352 686 -288
rect -686 -368 686 -352
rect -686 -432 602 -368
rect 666 -432 686 -368
rect -686 -448 686 -432
rect -686 -512 602 -448
rect 666 -512 686 -448
rect -686 -540 686 -512
<< via3 >>
rect 602 448 666 512
rect 602 368 666 432
rect 602 288 666 352
rect 602 208 666 272
rect 602 128 666 192
rect 602 48 666 112
rect 602 -32 666 32
rect 602 -112 666 -48
rect 602 -192 666 -128
rect 602 -272 666 -208
rect 602 -352 666 -288
rect 602 -432 666 -368
rect 602 -512 666 -448
<< mimcap >>
rect -646 432 354 500
rect -646 -432 -578 432
rect 286 -432 354 432
rect -646 -500 354 -432
<< mimcapcontact >>
rect -578 -432 286 432
<< metal4 >>
rect 586 512 682 528
rect -607 432 315 461
rect -607 -432 -578 432
rect 286 -432 315 432
rect -607 -461 315 -432
rect 586 448 602 512
rect 666 448 682 512
rect 586 432 682 448
rect 586 368 602 432
rect 666 368 682 432
rect 586 352 682 368
rect 586 288 602 352
rect 666 288 682 352
rect 586 272 682 288
rect 586 208 602 272
rect 666 208 682 272
rect 586 192 682 208
rect 586 128 602 192
rect 666 128 682 192
rect 586 112 682 128
rect 586 48 602 112
rect 666 48 682 112
rect 586 32 682 48
rect 586 -32 602 32
rect 666 -32 682 32
rect 586 -48 682 -32
rect 586 -112 602 -48
rect 666 -112 682 -48
rect 586 -128 682 -112
rect 586 -192 602 -128
rect 666 -192 682 -128
rect 586 -208 682 -192
rect 586 -272 602 -208
rect 666 -272 682 -208
rect 586 -288 682 -272
rect 586 -352 602 -288
rect 666 -352 682 -288
rect 586 -368 682 -352
rect 586 -432 602 -368
rect 666 -432 682 -368
rect 586 -448 682 -432
rect 586 -512 602 -448
rect 666 -512 682 -448
rect 586 -528 682 -512
<< properties >>
string FIXED_BBOX -686 -540 394 540
<< end >>
