magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< error_s >>
rect 12480 21853 12510 21951
rect 12226 21817 12625 21853
rect 12386 21783 12457 21817
rect 12423 21781 12457 21783
rect 12424 21377 12457 21781
rect 12460 21783 12648 21817
rect 12460 21747 12546 21783
rect 12460 21413 12493 21747
rect 12424 15163 12457 15166
rect 12460 15127 12493 15130
<< nwell >>
rect 367 21817 12422 21853
rect 12457 21817 12460 21853
rect 367 21413 12460 21817
rect 12480 21783 12510 21817
rect 367 21410 12493 21413
rect 367 20900 12500 21410
rect 367 20640 8190 20900
rect 9510 20640 12500 20900
rect 367 15130 12500 20640
rect 367 15127 12460 15130
<< pwell >>
rect 357 13157 11633 13243
rect 357 -657 443 13157
rect 2664 12230 2996 12430
rect 5564 12220 5896 12420
rect 11547 11043 11633 13157
rect 11547 10957 22523 11043
rect 14234 10314 14446 10466
rect 1564 5760 1716 5960
rect 1474 -657 1806 -410
rect 19114 -657 19266 -340
rect 21084 -657 21236 -350
rect 21454 -657 21606 -350
rect 22437 -657 22523 10957
rect 357 -743 22523 -657
<< psubdiff >>
rect 383 13183 458 13217
rect 492 13183 526 13217
rect 560 13183 594 13217
rect 628 13183 662 13217
rect 696 13183 730 13217
rect 764 13183 798 13217
rect 832 13183 866 13217
rect 900 13183 934 13217
rect 968 13183 1002 13217
rect 1036 13183 1070 13217
rect 1104 13183 1138 13217
rect 1172 13183 1206 13217
rect 1240 13183 1274 13217
rect 1308 13183 1342 13217
rect 1376 13183 1410 13217
rect 1444 13183 1478 13217
rect 1512 13183 1546 13217
rect 1580 13183 1614 13217
rect 1648 13183 1682 13217
rect 1716 13183 1750 13217
rect 1784 13183 1818 13217
rect 1852 13183 1886 13217
rect 1920 13183 1954 13217
rect 1988 13183 2022 13217
rect 2056 13183 2090 13217
rect 2124 13183 2158 13217
rect 2192 13183 2226 13217
rect 2260 13183 2294 13217
rect 2328 13183 2362 13217
rect 2396 13183 2430 13217
rect 2464 13183 2498 13217
rect 2532 13183 2566 13217
rect 2600 13183 2634 13217
rect 2668 13183 2702 13217
rect 2736 13183 2770 13217
rect 2804 13183 2838 13217
rect 2872 13183 2906 13217
rect 2940 13183 2974 13217
rect 3008 13183 3042 13217
rect 3076 13183 3110 13217
rect 3144 13183 3178 13217
rect 3212 13183 3246 13217
rect 3280 13183 3314 13217
rect 3348 13183 3382 13217
rect 3416 13183 3450 13217
rect 3484 13183 3518 13217
rect 3552 13183 3586 13217
rect 3620 13183 3654 13217
rect 3688 13183 3722 13217
rect 3756 13183 3790 13217
rect 3824 13183 3858 13217
rect 3892 13183 3926 13217
rect 3960 13183 3994 13217
rect 4028 13183 4062 13217
rect 4096 13183 4130 13217
rect 4164 13183 4198 13217
rect 4232 13183 4266 13217
rect 4300 13183 4334 13217
rect 4368 13183 4402 13217
rect 4436 13183 4470 13217
rect 4504 13183 4538 13217
rect 4572 13183 4606 13217
rect 4640 13183 4674 13217
rect 4708 13183 4742 13217
rect 4776 13183 4810 13217
rect 4844 13183 4878 13217
rect 4912 13183 4946 13217
rect 4980 13183 5014 13217
rect 5048 13183 5082 13217
rect 5116 13183 5150 13217
rect 5184 13183 5218 13217
rect 5252 13183 5286 13217
rect 5320 13183 5354 13217
rect 5388 13183 5422 13217
rect 5456 13183 5490 13217
rect 5524 13183 5558 13217
rect 5592 13183 5626 13217
rect 5660 13183 5694 13217
rect 5728 13183 5762 13217
rect 5796 13183 5830 13217
rect 5864 13183 5898 13217
rect 5932 13183 5966 13217
rect 6000 13183 6034 13217
rect 6068 13183 6102 13217
rect 6136 13183 6170 13217
rect 6204 13183 6238 13217
rect 6272 13183 6306 13217
rect 6340 13183 6374 13217
rect 6408 13183 6442 13217
rect 6476 13183 6510 13217
rect 6544 13183 6578 13217
rect 6612 13183 6646 13217
rect 6680 13183 6714 13217
rect 6748 13183 6782 13217
rect 6816 13183 6850 13217
rect 6884 13183 6918 13217
rect 6952 13183 6986 13217
rect 7020 13183 7054 13217
rect 7088 13183 7122 13217
rect 7156 13183 7190 13217
rect 7224 13183 7258 13217
rect 7292 13183 7326 13217
rect 7360 13183 7394 13217
rect 7428 13183 7462 13217
rect 7496 13183 7530 13217
rect 7564 13183 7598 13217
rect 7632 13183 7666 13217
rect 7700 13183 7734 13217
rect 7768 13183 7802 13217
rect 7836 13183 7870 13217
rect 7904 13183 7938 13217
rect 7972 13183 8006 13217
rect 8040 13183 8074 13217
rect 8108 13183 8142 13217
rect 8176 13183 8210 13217
rect 8244 13183 8278 13217
rect 8312 13183 8346 13217
rect 8380 13183 8414 13217
rect 8448 13183 8482 13217
rect 8516 13183 8550 13217
rect 8584 13183 8618 13217
rect 8652 13183 8686 13217
rect 8720 13183 8754 13217
rect 8788 13183 8822 13217
rect 8856 13183 8890 13217
rect 8924 13183 8958 13217
rect 8992 13183 9026 13217
rect 9060 13183 9094 13217
rect 9128 13183 9162 13217
rect 9196 13183 9230 13217
rect 9264 13183 9384 13217
rect 9418 13183 9452 13217
rect 9486 13183 9520 13217
rect 9554 13183 9588 13217
rect 9622 13183 9656 13217
rect 9690 13183 9724 13217
rect 9758 13183 9792 13217
rect 9826 13183 9860 13217
rect 9894 13183 9928 13217
rect 9962 13183 9996 13217
rect 10030 13183 10064 13217
rect 10098 13183 10132 13217
rect 10166 13183 10200 13217
rect 10234 13183 10268 13217
rect 10302 13183 10336 13217
rect 10370 13183 10404 13217
rect 10438 13183 10472 13217
rect 10506 13183 10540 13217
rect 10574 13183 10608 13217
rect 10642 13183 10676 13217
rect 10710 13183 10744 13217
rect 10778 13183 10812 13217
rect 10846 13183 10880 13217
rect 10914 13183 10948 13217
rect 10982 13183 11016 13217
rect 11050 13183 11084 13217
rect 11118 13183 11152 13217
rect 11186 13183 11220 13217
rect 11254 13183 11288 13217
rect 11322 13183 11356 13217
rect 11390 13183 11424 13217
rect 11458 13183 11492 13217
rect 11526 13183 11607 13217
rect 383 13135 417 13183
rect 383 13067 417 13101
rect 383 12999 417 13033
rect 383 12931 417 12965
rect 383 12863 417 12897
rect 383 12795 417 12829
rect 383 12727 417 12761
rect 383 12659 417 12693
rect 383 12591 417 12625
rect 383 12523 417 12557
rect 383 12455 417 12489
rect 383 12387 417 12421
rect 11573 13137 11607 13183
rect 11573 13069 11607 13103
rect 11573 13001 11607 13035
rect 11573 12933 11607 12967
rect 11573 12865 11607 12899
rect 11573 12797 11607 12831
rect 11573 12729 11607 12763
rect 11573 12661 11607 12695
rect 11573 12593 11607 12627
rect 11573 12525 11607 12559
rect 11573 12457 11607 12491
rect 383 12319 417 12353
rect 383 12251 417 12285
rect 2690 12347 2790 12404
rect 2690 12313 2723 12347
rect 2757 12313 2790 12347
rect 2690 12256 2790 12313
rect 2870 12347 2970 12404
rect 2870 12313 2903 12347
rect 2937 12313 2970 12347
rect 2870 12256 2970 12313
rect 5590 12337 5690 12394
rect 5590 12303 5623 12337
rect 5657 12303 5690 12337
rect 5590 12246 5690 12303
rect 5770 12337 5870 12394
rect 5770 12303 5803 12337
rect 5837 12303 5870 12337
rect 5770 12246 5870 12303
rect 11573 12389 11607 12423
rect 11573 12321 11607 12355
rect 11573 12253 11607 12287
rect 383 12183 417 12217
rect 383 12115 417 12149
rect 383 12047 417 12081
rect 383 11979 417 12013
rect 383 11911 417 11945
rect 383 11843 417 11877
rect 383 11775 417 11809
rect 383 11707 417 11741
rect 383 11639 417 11673
rect 383 11571 417 11605
rect 383 11503 417 11537
rect 383 11435 417 11469
rect 383 11367 417 11401
rect 383 11299 417 11333
rect 383 11231 417 11265
rect 383 11163 417 11197
rect 383 11095 417 11129
rect 383 11027 417 11061
rect 383 10959 417 10993
rect 11573 12185 11607 12219
rect 11573 12117 11607 12151
rect 11573 12049 11607 12083
rect 11573 11981 11607 12015
rect 11573 11913 11607 11947
rect 11573 11845 11607 11879
rect 11573 11777 11607 11811
rect 11573 11709 11607 11743
rect 11573 11641 11607 11675
rect 11573 11573 11607 11607
rect 11573 11505 11607 11539
rect 11573 11437 11607 11471
rect 11573 11369 11607 11403
rect 11573 11301 11607 11335
rect 11573 11233 11607 11267
rect 11573 11165 11607 11199
rect 11573 11097 11607 11131
rect 11573 11017 11607 11063
rect 11573 10983 11644 11017
rect 11678 10983 11712 11017
rect 11746 10983 11780 11017
rect 11814 10983 11848 11017
rect 11882 10983 11916 11017
rect 11950 10983 11984 11017
rect 12018 10983 12052 11017
rect 12086 10983 12120 11017
rect 12154 10983 12188 11017
rect 12222 10983 12256 11017
rect 12290 10983 12324 11017
rect 12358 10983 12392 11017
rect 12426 10983 12460 11017
rect 12494 10983 12528 11017
rect 12562 10983 12596 11017
rect 12630 10983 12664 11017
rect 12698 10983 12732 11017
rect 12766 10983 12800 11017
rect 12834 10983 12868 11017
rect 12902 10983 12936 11017
rect 12970 10983 13004 11017
rect 13038 10983 13072 11017
rect 13106 10983 13140 11017
rect 13174 10983 13208 11017
rect 13242 10983 13276 11017
rect 13310 10983 13344 11017
rect 13378 10983 13412 11017
rect 13446 10983 13480 11017
rect 13514 10983 13548 11017
rect 13582 10983 13616 11017
rect 13650 10983 13684 11017
rect 13718 10983 13752 11017
rect 13786 10983 13820 11017
rect 13854 10983 13888 11017
rect 13922 10983 13956 11017
rect 13990 10983 14024 11017
rect 14058 10983 14092 11017
rect 14126 10983 14160 11017
rect 14194 10983 14228 11017
rect 14262 10983 14296 11017
rect 14330 10983 14364 11017
rect 14398 10983 14432 11017
rect 14466 10983 14500 11017
rect 14534 10983 14568 11017
rect 14602 10983 14636 11017
rect 14670 10983 14704 11017
rect 14738 10983 14772 11017
rect 14806 10983 14840 11017
rect 14874 10983 14908 11017
rect 14942 10983 14976 11017
rect 15010 10983 15044 11017
rect 15078 10983 15112 11017
rect 15146 10983 15180 11017
rect 15214 10983 15248 11017
rect 15282 10983 15316 11017
rect 15350 10983 15384 11017
rect 15418 10983 15452 11017
rect 15486 10983 15520 11017
rect 15554 10983 15588 11017
rect 15622 10983 15656 11017
rect 15690 10983 15724 11017
rect 15758 10983 15792 11017
rect 15826 10983 15860 11017
rect 15894 10983 15928 11017
rect 15962 10983 15996 11017
rect 16030 10983 16064 11017
rect 16098 10983 16132 11017
rect 16166 10983 16200 11017
rect 16234 10983 16268 11017
rect 16302 10983 16336 11017
rect 16370 10983 16404 11017
rect 16438 10983 16472 11017
rect 16506 10983 16540 11017
rect 16574 10983 16608 11017
rect 16642 10983 16676 11017
rect 16710 10983 16744 11017
rect 16778 10983 16812 11017
rect 16846 10983 16880 11017
rect 16914 10983 16948 11017
rect 16982 10983 17016 11017
rect 17050 10983 17084 11017
rect 17118 10983 17152 11017
rect 17186 10983 17220 11017
rect 17254 10983 17288 11017
rect 17322 10983 17356 11017
rect 17390 10983 17424 11017
rect 17458 10983 17492 11017
rect 17526 10983 17560 11017
rect 17594 10983 17628 11017
rect 17662 10983 17696 11017
rect 17730 10983 17764 11017
rect 17798 10983 17832 11017
rect 17866 10983 17900 11017
rect 17934 10983 17968 11017
rect 18002 10983 18036 11017
rect 18070 10983 18104 11017
rect 18138 10983 18172 11017
rect 18206 10983 18240 11017
rect 18274 10983 18308 11017
rect 18342 10983 18376 11017
rect 18410 10983 18444 11017
rect 18478 10983 18512 11017
rect 18546 10983 18580 11017
rect 18614 10983 18648 11017
rect 18682 10983 18716 11017
rect 18750 10983 18784 11017
rect 18818 10983 18852 11017
rect 18886 10983 18920 11017
rect 18954 10983 18988 11017
rect 19022 10983 19056 11017
rect 19090 10983 19124 11017
rect 19158 10983 19192 11017
rect 19226 10983 19260 11017
rect 19294 10983 19328 11017
rect 19362 10983 19396 11017
rect 19430 10983 19464 11017
rect 19498 10983 19532 11017
rect 19566 10983 19600 11017
rect 19634 10983 19668 11017
rect 19702 10983 19736 11017
rect 19770 10983 19804 11017
rect 19838 10983 19872 11017
rect 19906 10983 19940 11017
rect 19974 10983 20008 11017
rect 20042 10983 20076 11017
rect 20110 10983 20144 11017
rect 20178 10983 20212 11017
rect 20246 10983 20280 11017
rect 20314 10983 20348 11017
rect 20382 10983 20416 11017
rect 20450 10983 20484 11017
rect 20518 10983 20552 11017
rect 20586 10983 20620 11017
rect 20654 10983 20688 11017
rect 20722 10983 20756 11017
rect 20790 10983 20824 11017
rect 20858 10983 20892 11017
rect 20926 10983 20960 11017
rect 20994 10983 21028 11017
rect 21062 10983 21096 11017
rect 21130 10983 21164 11017
rect 21198 10983 21232 11017
rect 21266 10983 21300 11017
rect 21334 10983 21368 11017
rect 21402 10983 21436 11017
rect 21470 10983 21504 11017
rect 21538 10983 21572 11017
rect 21606 10983 21640 11017
rect 21674 10983 21708 11017
rect 21742 10983 21776 11017
rect 21810 10983 21844 11017
rect 21878 10983 21912 11017
rect 21946 10983 21980 11017
rect 22014 10983 22048 11017
rect 22082 10983 22116 11017
rect 22150 10983 22184 11017
rect 22218 10983 22252 11017
rect 22286 10983 22320 11017
rect 22354 10983 22388 11017
rect 22422 10983 22497 11017
rect 383 10891 417 10925
rect 383 10823 417 10857
rect 383 10755 417 10789
rect 383 10687 417 10721
rect 383 10619 417 10653
rect 383 10551 417 10585
rect 383 10483 417 10517
rect 383 10415 417 10449
rect 22463 10947 22497 10983
rect 22463 10879 22497 10913
rect 22463 10811 22497 10845
rect 22463 10743 22497 10777
rect 22463 10675 22497 10709
rect 22463 10607 22497 10641
rect 22463 10539 22497 10573
rect 22463 10471 22497 10505
rect 383 10347 417 10381
rect 14260 10407 14420 10440
rect 14260 10373 14323 10407
rect 14357 10373 14420 10407
rect 14260 10340 14420 10373
rect 22463 10403 22497 10437
rect 383 10279 417 10313
rect 383 10211 417 10245
rect 383 10143 417 10177
rect 383 10075 417 10109
rect 383 10007 417 10041
rect 383 9939 417 9973
rect 383 9871 417 9905
rect 383 9803 417 9837
rect 383 9735 417 9769
rect 383 9667 417 9701
rect 383 9599 417 9633
rect 383 9531 417 9565
rect 383 9463 417 9497
rect 383 9395 417 9429
rect 383 9327 417 9361
rect 383 9259 417 9293
rect 383 9191 417 9225
rect 383 9123 417 9157
rect 383 9055 417 9089
rect 383 8987 417 9021
rect 383 8919 417 8953
rect 383 8851 417 8885
rect 383 8783 417 8817
rect 383 8715 417 8749
rect 383 8647 417 8681
rect 383 8579 417 8613
rect 383 8511 417 8545
rect 383 8443 417 8477
rect 383 8375 417 8409
rect 383 8307 417 8341
rect 383 8239 417 8273
rect 383 8171 417 8205
rect 383 8103 417 8137
rect 383 8035 417 8069
rect 383 7967 417 8001
rect 383 7899 417 7933
rect 383 7831 417 7865
rect 383 7763 417 7797
rect 383 7695 417 7729
rect 383 7627 417 7661
rect 383 7559 417 7593
rect 383 7491 417 7525
rect 383 7423 417 7457
rect 383 7355 417 7389
rect 383 7287 417 7321
rect 383 7219 417 7253
rect 383 7151 417 7185
rect 383 7083 417 7117
rect 383 7015 417 7049
rect 383 6947 417 6981
rect 383 6879 417 6913
rect 383 6811 417 6845
rect 383 6743 417 6777
rect 383 6675 417 6709
rect 383 6607 417 6641
rect 383 6539 417 6573
rect 383 6471 417 6505
rect 383 6403 417 6437
rect 383 6335 417 6369
rect 383 6267 417 6301
rect 383 6199 417 6233
rect 383 6131 417 6165
rect 383 6063 417 6097
rect 383 5995 417 6029
rect 383 5927 417 5961
rect 22463 10335 22497 10369
rect 22463 10267 22497 10301
rect 22463 10199 22497 10233
rect 22463 10131 22497 10165
rect 22463 10063 22497 10097
rect 22463 9995 22497 10029
rect 22463 9927 22497 9961
rect 22463 9859 22497 9893
rect 22463 9791 22497 9825
rect 22463 9723 22497 9757
rect 22463 9655 22497 9689
rect 22463 9587 22497 9621
rect 22463 9519 22497 9553
rect 22463 9451 22497 9485
rect 22463 9383 22497 9417
rect 22463 9315 22497 9349
rect 22463 9247 22497 9281
rect 22463 9179 22497 9213
rect 22463 9111 22497 9145
rect 22463 9043 22497 9077
rect 22463 8975 22497 9009
rect 22463 8907 22497 8941
rect 22463 8839 22497 8873
rect 22463 8771 22497 8805
rect 22463 8703 22497 8737
rect 22463 8635 22497 8669
rect 22463 8567 22497 8601
rect 22463 8499 22497 8533
rect 22463 8431 22497 8465
rect 22463 8363 22497 8397
rect 22463 8295 22497 8329
rect 22463 8227 22497 8261
rect 22463 8159 22497 8193
rect 22463 8091 22497 8125
rect 22463 8023 22497 8057
rect 22463 7955 22497 7989
rect 22463 7887 22497 7921
rect 22463 7819 22497 7853
rect 22463 7751 22497 7785
rect 22463 7683 22497 7717
rect 22463 7615 22497 7649
rect 22463 7547 22497 7581
rect 22463 7479 22497 7513
rect 22463 7411 22497 7445
rect 22463 7343 22497 7377
rect 22463 7275 22497 7309
rect 22463 7207 22497 7241
rect 22463 7139 22497 7173
rect 22463 7071 22497 7105
rect 22463 7003 22497 7037
rect 22463 6935 22497 6969
rect 22463 6867 22497 6901
rect 22463 6799 22497 6833
rect 22463 6731 22497 6765
rect 22463 6663 22497 6697
rect 22463 6595 22497 6629
rect 22463 6527 22497 6561
rect 22463 6459 22497 6493
rect 22463 6391 22497 6425
rect 22463 6323 22497 6357
rect 22463 6255 22497 6289
rect 22463 6187 22497 6221
rect 22463 6119 22497 6153
rect 22463 6051 22497 6085
rect 22463 5983 22497 6017
rect 383 5859 417 5893
rect 383 5791 417 5825
rect 1590 5877 1690 5934
rect 1590 5843 1623 5877
rect 1657 5843 1690 5877
rect 1590 5786 1690 5843
rect 22463 5915 22497 5949
rect 22463 5847 22497 5881
rect 383 5723 417 5757
rect 383 5655 417 5689
rect 383 5587 417 5621
rect 383 5519 417 5553
rect 383 5451 417 5485
rect 383 5383 417 5417
rect 383 5315 417 5349
rect 383 5247 417 5281
rect 383 5179 417 5213
rect 383 5111 417 5145
rect 383 5043 417 5077
rect 383 4975 417 5009
rect 383 4907 417 4941
rect 383 4839 417 4873
rect 383 4771 417 4805
rect 383 4703 417 4737
rect 383 4635 417 4669
rect 383 4567 417 4601
rect 383 4499 417 4533
rect 383 4431 417 4465
rect 383 4363 417 4397
rect 383 4295 417 4329
rect 383 4227 417 4261
rect 383 4159 417 4193
rect 383 4091 417 4125
rect 383 4023 417 4057
rect 383 3955 417 3989
rect 383 3887 417 3921
rect 383 3819 417 3853
rect 383 3751 417 3785
rect 383 3683 417 3717
rect 383 3615 417 3649
rect 383 3547 417 3581
rect 383 3479 417 3513
rect 383 3411 417 3445
rect 383 3343 417 3377
rect 383 3275 417 3309
rect 383 3207 417 3241
rect 383 3139 417 3173
rect 383 3071 417 3105
rect 383 3003 417 3037
rect 383 2935 417 2969
rect 383 2867 417 2901
rect 383 2799 417 2833
rect 383 2731 417 2765
rect 383 2663 417 2697
rect 383 2595 417 2629
rect 383 2527 417 2561
rect 383 2459 417 2493
rect 383 2391 417 2425
rect 383 2323 417 2357
rect 383 2255 417 2289
rect 383 2187 417 2221
rect 383 2119 417 2153
rect 383 2051 417 2085
rect 383 1983 417 2017
rect 383 1915 417 1949
rect 383 1847 417 1881
rect 383 1779 417 1813
rect 383 1711 417 1745
rect 383 1643 417 1677
rect 383 1575 417 1609
rect 383 1507 417 1541
rect 383 1439 417 1473
rect 383 1371 417 1405
rect 383 1303 417 1337
rect 383 1235 417 1269
rect 383 1167 417 1201
rect 383 1099 417 1133
rect 383 1031 417 1065
rect 383 963 417 997
rect 383 895 417 929
rect 383 827 417 861
rect 383 759 417 793
rect 383 691 417 725
rect 383 623 417 657
rect 383 555 417 589
rect 383 487 417 521
rect 383 419 417 453
rect 383 351 417 385
rect 383 283 417 317
rect 383 215 417 249
rect 383 147 417 181
rect 383 79 417 113
rect 383 11 417 45
rect 383 -57 417 -23
rect 383 -125 417 -91
rect 383 -193 417 -159
rect 383 -261 417 -227
rect 383 -329 417 -295
rect 383 -397 417 -363
rect 22463 5779 22497 5813
rect 22463 5711 22497 5745
rect 22463 5643 22497 5677
rect 22463 5575 22497 5609
rect 22463 5507 22497 5541
rect 22463 5439 22497 5473
rect 22463 5371 22497 5405
rect 22463 5303 22497 5337
rect 22463 5235 22497 5269
rect 22463 5167 22497 5201
rect 22463 5099 22497 5133
rect 22463 5031 22497 5065
rect 22463 4963 22497 4997
rect 22463 4895 22497 4929
rect 22463 4827 22497 4861
rect 22463 4759 22497 4793
rect 22463 4691 22497 4725
rect 22463 4623 22497 4657
rect 22463 4555 22497 4589
rect 22463 4487 22497 4521
rect 22463 4419 22497 4453
rect 22463 4351 22497 4385
rect 22463 4283 22497 4317
rect 22463 4215 22497 4249
rect 22463 4147 22497 4181
rect 22463 4079 22497 4113
rect 22463 4011 22497 4045
rect 22463 3943 22497 3977
rect 22463 3875 22497 3909
rect 22463 3807 22497 3841
rect 22463 3739 22497 3773
rect 22463 3671 22497 3705
rect 22463 3603 22497 3637
rect 22463 3535 22497 3569
rect 22463 3467 22497 3501
rect 22463 3399 22497 3433
rect 22463 3331 22497 3365
rect 22463 3263 22497 3297
rect 22463 3195 22497 3229
rect 22463 3127 22497 3161
rect 22463 3059 22497 3093
rect 22463 2991 22497 3025
rect 22463 2923 22497 2957
rect 22463 2855 22497 2889
rect 22463 2787 22497 2821
rect 22463 2719 22497 2753
rect 22463 2651 22497 2685
rect 22463 2583 22497 2617
rect 22463 2515 22497 2549
rect 22463 2447 22497 2481
rect 22463 2379 22497 2413
rect 22463 2311 22497 2345
rect 22463 2243 22497 2277
rect 22463 2175 22497 2209
rect 22463 2107 22497 2141
rect 22463 2039 22497 2073
rect 22463 1971 22497 2005
rect 22463 1903 22497 1937
rect 22463 1835 22497 1869
rect 22463 1767 22497 1801
rect 22463 1699 22497 1733
rect 22463 1631 22497 1665
rect 22463 1563 22497 1597
rect 22463 1495 22497 1529
rect 22463 1427 22497 1461
rect 22463 1359 22497 1393
rect 22463 1291 22497 1325
rect 22463 1223 22497 1257
rect 22463 1155 22497 1189
rect 22463 1087 22497 1121
rect 22463 1019 22497 1053
rect 22463 951 22497 985
rect 22463 883 22497 917
rect 22463 815 22497 849
rect 22463 747 22497 781
rect 22463 679 22497 713
rect 22463 611 22497 645
rect 22463 543 22497 577
rect 22463 475 22497 509
rect 22463 407 22497 441
rect 22463 339 22497 373
rect 22463 271 22497 305
rect 22463 203 22497 237
rect 22463 135 22497 169
rect 22463 67 22497 101
rect 22463 -1 22497 33
rect 22463 -69 22497 -35
rect 22463 -137 22497 -103
rect 22463 -205 22497 -171
rect 22463 -273 22497 -239
rect 22463 -341 22497 -307
rect 383 -465 417 -431
rect 19140 -423 19240 -366
rect 383 -533 417 -499
rect 383 -601 417 -567
rect 1500 -493 1600 -436
rect 1500 -527 1533 -493
rect 1567 -527 1600 -493
rect 1500 -584 1600 -527
rect 1680 -493 1780 -436
rect 1680 -527 1713 -493
rect 1747 -527 1780 -493
rect 19140 -457 19173 -423
rect 19207 -457 19240 -423
rect 19140 -514 19240 -457
rect 21110 -433 21210 -376
rect 21110 -467 21143 -433
rect 21177 -467 21210 -433
rect 21110 -524 21210 -467
rect 21480 -433 21580 -376
rect 21480 -467 21513 -433
rect 21547 -467 21580 -433
rect 21480 -524 21580 -467
rect 22463 -409 22497 -375
rect 22463 -477 22497 -443
rect 1680 -584 1780 -527
rect 22463 -545 22497 -511
rect 383 -683 417 -635
rect 22463 -613 22497 -579
rect 22463 -683 22497 -647
rect 383 -717 475 -683
rect 509 -717 543 -683
rect 577 -717 611 -683
rect 645 -717 679 -683
rect 713 -717 747 -683
rect 781 -717 815 -683
rect 849 -717 883 -683
rect 917 -717 951 -683
rect 985 -717 1019 -683
rect 1053 -717 1087 -683
rect 1121 -717 1155 -683
rect 1189 -717 1223 -683
rect 1257 -717 1291 -683
rect 1325 -717 1359 -683
rect 1393 -717 1427 -683
rect 1461 -717 1495 -683
rect 1529 -717 1563 -683
rect 1597 -717 1631 -683
rect 1665 -717 1699 -683
rect 1733 -717 1767 -683
rect 1801 -717 1835 -683
rect 1869 -717 1903 -683
rect 1937 -717 1971 -683
rect 2005 -717 2039 -683
rect 2073 -717 2107 -683
rect 2141 -717 2175 -683
rect 2209 -717 2243 -683
rect 2277 -717 2311 -683
rect 2345 -717 2379 -683
rect 2413 -717 2447 -683
rect 2481 -717 2515 -683
rect 2549 -717 2583 -683
rect 2617 -717 2651 -683
rect 2685 -717 2719 -683
rect 2753 -717 2787 -683
rect 2821 -717 2855 -683
rect 2889 -717 2923 -683
rect 2957 -717 2991 -683
rect 3025 -717 3059 -683
rect 3093 -717 3127 -683
rect 3161 -717 3195 -683
rect 3229 -717 3263 -683
rect 3297 -717 3331 -683
rect 3365 -717 3399 -683
rect 3433 -717 3467 -683
rect 3501 -717 3535 -683
rect 3569 -717 3603 -683
rect 3637 -717 3671 -683
rect 3705 -717 3739 -683
rect 3773 -717 3807 -683
rect 3841 -717 3875 -683
rect 3909 -717 3943 -683
rect 3977 -717 4011 -683
rect 4045 -717 4079 -683
rect 4113 -717 4147 -683
rect 4181 -717 4215 -683
rect 4249 -717 4283 -683
rect 4317 -717 4351 -683
rect 4385 -717 4419 -683
rect 4453 -717 4487 -683
rect 4521 -717 4555 -683
rect 4589 -717 4623 -683
rect 4657 -717 4691 -683
rect 4725 -717 4759 -683
rect 4793 -717 4827 -683
rect 4861 -717 4895 -683
rect 4929 -717 4963 -683
rect 4997 -717 5031 -683
rect 5065 -717 5099 -683
rect 5133 -717 5167 -683
rect 5201 -717 5235 -683
rect 5269 -717 5303 -683
rect 5337 -717 5371 -683
rect 5405 -717 5439 -683
rect 5473 -717 5507 -683
rect 5541 -717 5575 -683
rect 5609 -717 5643 -683
rect 5677 -717 5711 -683
rect 5745 -717 5779 -683
rect 5813 -717 5847 -683
rect 5881 -717 5915 -683
rect 5949 -717 5983 -683
rect 6017 -717 6051 -683
rect 6085 -717 6119 -683
rect 6153 -717 6187 -683
rect 6221 -717 6255 -683
rect 6289 -717 6323 -683
rect 6357 -717 6391 -683
rect 6425 -717 6459 -683
rect 6493 -717 6527 -683
rect 6561 -717 6595 -683
rect 6629 -717 6663 -683
rect 6697 -717 6731 -683
rect 6765 -717 6799 -683
rect 6833 -717 6867 -683
rect 6901 -717 6935 -683
rect 6969 -717 7003 -683
rect 7037 -717 7071 -683
rect 7105 -717 7139 -683
rect 7173 -717 7207 -683
rect 7241 -717 7275 -683
rect 7309 -717 7343 -683
rect 7377 -717 7411 -683
rect 7445 -717 7479 -683
rect 7513 -717 7547 -683
rect 7581 -717 7615 -683
rect 7649 -717 7683 -683
rect 7717 -717 7751 -683
rect 7785 -717 7819 -683
rect 7853 -717 7887 -683
rect 7921 -717 7955 -683
rect 7989 -717 8023 -683
rect 8057 -717 8091 -683
rect 8125 -717 8159 -683
rect 8193 -717 8227 -683
rect 8261 -717 8295 -683
rect 8329 -717 8363 -683
rect 8397 -717 8431 -683
rect 8465 -717 8499 -683
rect 8533 -717 8567 -683
rect 8601 -717 8635 -683
rect 8669 -717 8703 -683
rect 8737 -717 8771 -683
rect 8805 -717 8839 -683
rect 8873 -717 8907 -683
rect 8941 -717 8975 -683
rect 9009 -717 9043 -683
rect 9077 -717 9111 -683
rect 9145 -717 9179 -683
rect 9213 -717 9247 -683
rect 9281 -717 9315 -683
rect 9349 -717 9383 -683
rect 9417 -717 9451 -683
rect 9485 -717 9519 -683
rect 9553 -717 9587 -683
rect 9621 -717 9655 -683
rect 9689 -717 9723 -683
rect 9757 -717 9791 -683
rect 9825 -717 9859 -683
rect 9893 -717 9927 -683
rect 9961 -717 9995 -683
rect 10029 -717 10063 -683
rect 10097 -717 10131 -683
rect 10165 -717 10199 -683
rect 10233 -717 10267 -683
rect 10301 -717 10335 -683
rect 10369 -717 10403 -683
rect 10437 -717 10471 -683
rect 10505 -717 10539 -683
rect 10573 -717 10607 -683
rect 10641 -717 10675 -683
rect 10709 -717 10743 -683
rect 10777 -717 10811 -683
rect 10845 -717 10879 -683
rect 10913 -717 10947 -683
rect 10981 -717 11015 -683
rect 11049 -717 11083 -683
rect 11117 -717 11151 -683
rect 11185 -717 11219 -683
rect 11253 -717 11287 -683
rect 11321 -717 11355 -683
rect 11389 -717 11423 -683
rect 11457 -717 11491 -683
rect 11525 -717 11559 -683
rect 11593 -717 11627 -683
rect 11661 -717 11695 -683
rect 11729 -717 11763 -683
rect 11797 -717 11831 -683
rect 11865 -717 11899 -683
rect 11933 -717 11967 -683
rect 12001 -717 12035 -683
rect 12069 -717 12103 -683
rect 12137 -717 12171 -683
rect 12205 -717 12239 -683
rect 12273 -717 12307 -683
rect 12341 -717 12375 -683
rect 12409 -717 12443 -683
rect 12477 -717 12511 -683
rect 12545 -717 12579 -683
rect 12613 -717 12647 -683
rect 12681 -717 12715 -683
rect 12749 -717 12783 -683
rect 12817 -717 12851 -683
rect 12885 -717 12919 -683
rect 12953 -717 12987 -683
rect 13021 -717 13055 -683
rect 13089 -717 13123 -683
rect 13157 -717 13191 -683
rect 13225 -717 13259 -683
rect 13293 -717 13327 -683
rect 13361 -717 13395 -683
rect 13429 -717 13463 -683
rect 13497 -717 13531 -683
rect 13565 -717 13599 -683
rect 13633 -717 13667 -683
rect 13701 -717 13735 -683
rect 13769 -717 13803 -683
rect 13837 -717 13871 -683
rect 13905 -717 13939 -683
rect 13973 -717 14007 -683
rect 14041 -717 14075 -683
rect 14109 -717 14143 -683
rect 14177 -717 14211 -683
rect 14245 -717 14279 -683
rect 14313 -717 14347 -683
rect 14381 -717 14415 -683
rect 14449 -717 14483 -683
rect 14517 -717 14551 -683
rect 14585 -717 14619 -683
rect 14653 -717 14687 -683
rect 14721 -717 14755 -683
rect 14789 -717 14823 -683
rect 14857 -717 14891 -683
rect 14925 -717 14959 -683
rect 14993 -717 15027 -683
rect 15061 -717 15095 -683
rect 15129 -717 15163 -683
rect 15197 -717 15231 -683
rect 15265 -717 15299 -683
rect 15333 -717 15367 -683
rect 15401 -717 15435 -683
rect 15469 -717 15503 -683
rect 15537 -717 15571 -683
rect 15605 -717 15639 -683
rect 15673 -717 15707 -683
rect 15741 -717 15775 -683
rect 15809 -717 15843 -683
rect 15877 -717 15911 -683
rect 15945 -717 15979 -683
rect 16013 -717 16047 -683
rect 16081 -717 16115 -683
rect 16149 -717 16183 -683
rect 16217 -717 16251 -683
rect 16285 -717 16319 -683
rect 16353 -717 16387 -683
rect 16421 -717 16455 -683
rect 16489 -717 16523 -683
rect 16557 -717 16591 -683
rect 16625 -717 16659 -683
rect 16693 -717 16727 -683
rect 16761 -717 16795 -683
rect 16829 -717 16863 -683
rect 16897 -717 16931 -683
rect 16965 -717 16999 -683
rect 17033 -717 17067 -683
rect 17101 -717 17135 -683
rect 17169 -717 17203 -683
rect 17237 -717 17271 -683
rect 17305 -717 17339 -683
rect 17373 -717 17407 -683
rect 17441 -717 17475 -683
rect 17509 -717 17543 -683
rect 17577 -717 17611 -683
rect 17645 -717 17679 -683
rect 17713 -717 17747 -683
rect 17781 -717 17815 -683
rect 17849 -717 17883 -683
rect 17917 -717 17951 -683
rect 17985 -717 18019 -683
rect 18053 -717 18087 -683
rect 18121 -717 18155 -683
rect 18189 -717 18223 -683
rect 18257 -717 18291 -683
rect 18325 -717 18359 -683
rect 18393 -717 18427 -683
rect 18461 -717 18495 -683
rect 18529 -717 18563 -683
rect 18597 -717 18631 -683
rect 18665 -717 18699 -683
rect 18733 -717 18767 -683
rect 18801 -717 18835 -683
rect 18869 -717 18903 -683
rect 18937 -717 18971 -683
rect 19005 -717 19039 -683
rect 19073 -717 19107 -683
rect 19141 -717 19175 -683
rect 19209 -717 19243 -683
rect 19277 -717 19311 -683
rect 19345 -717 19379 -683
rect 19413 -717 19447 -683
rect 19481 -717 19515 -683
rect 19549 -717 19583 -683
rect 19617 -717 19651 -683
rect 19685 -717 19719 -683
rect 19753 -717 19787 -683
rect 19821 -717 19855 -683
rect 19889 -717 19923 -683
rect 19957 -717 19991 -683
rect 20025 -717 20059 -683
rect 20093 -717 20127 -683
rect 20161 -717 20195 -683
rect 20229 -717 20263 -683
rect 20297 -717 20331 -683
rect 20365 -717 20399 -683
rect 20433 -717 20467 -683
rect 20501 -717 20535 -683
rect 20569 -717 20603 -683
rect 20637 -717 20671 -683
rect 20705 -717 20739 -683
rect 20773 -717 20807 -683
rect 20841 -717 20875 -683
rect 20909 -717 20943 -683
rect 20977 -717 21011 -683
rect 21045 -717 21079 -683
rect 21113 -717 21147 -683
rect 21181 -717 21215 -683
rect 21249 -717 21283 -683
rect 21317 -717 21351 -683
rect 21385 -717 21419 -683
rect 21453 -717 21487 -683
rect 21521 -717 21555 -683
rect 21589 -717 21623 -683
rect 21657 -717 21691 -683
rect 21725 -717 21759 -683
rect 21793 -717 21827 -683
rect 21861 -717 21895 -683
rect 21929 -717 21963 -683
rect 21997 -717 22031 -683
rect 22065 -717 22099 -683
rect 22133 -717 22167 -683
rect 22201 -717 22235 -683
rect 22269 -717 22303 -683
rect 22337 -717 22371 -683
rect 22405 -717 22497 -683
<< nsubdiff >>
rect 403 21787 540 21817
rect 437 21783 540 21787
rect 574 21783 608 21817
rect 642 21783 676 21817
rect 710 21783 744 21817
rect 778 21783 812 21817
rect 846 21783 880 21817
rect 914 21783 948 21817
rect 982 21783 1016 21817
rect 1050 21783 1084 21817
rect 1118 21783 1152 21817
rect 1186 21783 1220 21817
rect 1254 21783 1288 21817
rect 1322 21783 1356 21817
rect 1390 21783 1424 21817
rect 1458 21783 1492 21817
rect 1526 21783 1560 21817
rect 1594 21783 1628 21817
rect 1662 21783 1696 21817
rect 1730 21783 1764 21817
rect 1798 21783 1832 21817
rect 1866 21783 1900 21817
rect 1934 21783 1968 21817
rect 2002 21783 2036 21817
rect 2070 21783 2104 21817
rect 2138 21783 2172 21817
rect 2206 21783 2240 21817
rect 2274 21783 2308 21817
rect 2342 21783 2376 21817
rect 2410 21783 2444 21817
rect 2478 21783 2512 21817
rect 2546 21783 2580 21817
rect 2614 21783 2648 21817
rect 2682 21783 2716 21817
rect 2750 21783 2784 21817
rect 2818 21783 2852 21817
rect 2886 21783 2920 21817
rect 2954 21783 2988 21817
rect 3022 21783 3056 21817
rect 3090 21783 3124 21817
rect 3158 21783 3192 21817
rect 3226 21783 3260 21817
rect 3294 21783 3328 21817
rect 3362 21783 3396 21817
rect 3430 21783 3464 21817
rect 3498 21783 3532 21817
rect 3566 21783 3600 21817
rect 3634 21783 3668 21817
rect 3702 21783 3736 21817
rect 3770 21783 3804 21817
rect 3838 21783 3872 21817
rect 3906 21783 3940 21817
rect 3974 21783 4008 21817
rect 4042 21783 4076 21817
rect 4110 21783 4144 21817
rect 4178 21783 4212 21817
rect 4246 21783 4280 21817
rect 4314 21783 4348 21817
rect 4382 21783 4416 21817
rect 4450 21783 4484 21817
rect 4518 21783 4552 21817
rect 4586 21783 4620 21817
rect 4654 21783 4688 21817
rect 4722 21783 4756 21817
rect 4790 21783 4824 21817
rect 4858 21783 4892 21817
rect 4926 21783 4960 21817
rect 4994 21783 5028 21817
rect 5062 21783 5096 21817
rect 5130 21783 5164 21817
rect 5198 21783 5232 21817
rect 5266 21783 5300 21817
rect 5334 21783 5368 21817
rect 5402 21783 5436 21817
rect 5470 21783 5504 21817
rect 5538 21783 5572 21817
rect 5606 21783 5640 21817
rect 5674 21783 5708 21817
rect 5742 21783 5776 21817
rect 5810 21783 5844 21817
rect 5878 21783 5912 21817
rect 5946 21783 5980 21817
rect 6014 21783 6048 21817
rect 6082 21783 6116 21817
rect 6150 21783 6184 21817
rect 6218 21783 6252 21817
rect 6286 21783 6320 21817
rect 6354 21783 6388 21817
rect 6422 21783 6456 21817
rect 6490 21783 6524 21817
rect 6558 21783 6592 21817
rect 6626 21783 6660 21817
rect 6694 21783 6728 21817
rect 6762 21783 6796 21817
rect 6830 21783 6864 21817
rect 6898 21783 6932 21817
rect 6966 21783 7000 21817
rect 7034 21783 7068 21817
rect 7102 21783 7136 21817
rect 7170 21783 7204 21817
rect 7238 21783 7272 21817
rect 7306 21783 7340 21817
rect 7374 21783 7408 21817
rect 7442 21783 7476 21817
rect 7510 21783 7544 21817
rect 7578 21783 7612 21817
rect 7646 21783 7680 21817
rect 7714 21783 7748 21817
rect 7782 21783 7816 21817
rect 7850 21783 7884 21817
rect 7918 21783 7952 21817
rect 7986 21783 8020 21817
rect 8054 21783 8088 21817
rect 8122 21783 8156 21817
rect 8190 21783 8224 21817
rect 8258 21783 8292 21817
rect 8326 21783 8360 21817
rect 8394 21783 8428 21817
rect 8462 21783 8496 21817
rect 8530 21783 8564 21817
rect 8598 21783 8632 21817
rect 8666 21783 8700 21817
rect 8734 21783 8768 21817
rect 8802 21783 8836 21817
rect 8870 21783 8904 21817
rect 8938 21783 8972 21817
rect 9006 21783 9040 21817
rect 9074 21783 9108 21817
rect 9142 21783 9176 21817
rect 9210 21783 9244 21817
rect 9278 21783 9312 21817
rect 9346 21783 9380 21817
rect 9414 21783 9448 21817
rect 9482 21783 9516 21817
rect 9550 21783 9584 21817
rect 9618 21783 9652 21817
rect 9686 21783 9720 21817
rect 9754 21783 9788 21817
rect 9822 21783 9856 21817
rect 9890 21783 9924 21817
rect 9958 21783 9992 21817
rect 10026 21783 10060 21817
rect 10094 21783 10128 21817
rect 10162 21783 10196 21817
rect 10230 21783 10264 21817
rect 10298 21783 10332 21817
rect 10366 21783 10400 21817
rect 10434 21783 10468 21817
rect 10502 21783 10536 21817
rect 10570 21783 10604 21817
rect 10638 21783 10672 21817
rect 10706 21783 10740 21817
rect 10774 21783 10808 21817
rect 10842 21783 10876 21817
rect 10910 21783 10944 21817
rect 10978 21783 11012 21817
rect 11046 21783 11080 21817
rect 11114 21783 11148 21817
rect 11182 21783 11216 21817
rect 11250 21783 11284 21817
rect 11318 21783 11352 21817
rect 11386 21783 11420 21817
rect 11454 21783 11488 21817
rect 11522 21783 11556 21817
rect 11590 21783 11624 21817
rect 11658 21783 11692 21817
rect 11726 21783 11760 21817
rect 11794 21783 11828 21817
rect 11862 21783 11896 21817
rect 11930 21783 11964 21817
rect 11998 21783 12032 21817
rect 12066 21783 12100 21817
rect 12134 21783 12168 21817
rect 12202 21783 12236 21817
rect 12270 21783 12304 21817
rect 12338 21783 12457 21817
rect 12480 21783 12510 21817
rect 403 21719 437 21753
rect 403 21651 437 21685
rect 403 21583 437 21617
rect 403 21515 437 21549
rect 403 21447 437 21481
rect 12423 21733 12457 21783
rect 12423 21665 12457 21699
rect 12423 21597 12457 21631
rect 12423 21529 12457 21563
rect 403 21379 437 21413
rect 1030 21442 1280 21470
rect 1030 21408 1075 21442
rect 1109 21408 1143 21442
rect 1177 21408 1211 21442
rect 1245 21408 1280 21442
rect 1030 21380 1280 21408
rect 7010 21437 7280 21470
rect 7010 21403 7055 21437
rect 7089 21403 7123 21437
rect 7157 21403 7191 21437
rect 7225 21403 7280 21437
rect 7010 21370 7280 21403
rect 12423 21461 12457 21495
rect 12423 21393 12457 21427
rect 403 21311 437 21345
rect 403 21243 437 21277
rect 403 21175 437 21209
rect 403 21107 437 21141
rect 403 21039 437 21073
rect 403 20971 437 21005
rect 403 20903 437 20937
rect 403 20835 437 20869
rect 403 20767 437 20801
rect 403 20699 437 20733
rect 403 20631 437 20665
rect 403 20563 437 20597
rect 403 20495 437 20529
rect 403 20427 437 20461
rect 403 20359 437 20393
rect 403 20291 437 20325
rect 403 20223 437 20257
rect 403 20155 437 20189
rect 403 20087 437 20121
rect 403 20019 437 20053
rect 403 19951 437 19985
rect 403 19883 437 19917
rect 403 19815 437 19849
rect 403 19747 437 19781
rect 403 19679 437 19713
rect 403 19611 437 19645
rect 403 19543 437 19577
rect 403 19475 437 19509
rect 403 19407 437 19441
rect 403 19339 437 19373
rect 403 19271 437 19305
rect 403 19203 437 19237
rect 403 19135 437 19169
rect 403 19067 437 19101
rect 403 18999 437 19033
rect 403 18931 437 18965
rect 403 18863 437 18897
rect 403 18795 437 18829
rect 403 18727 437 18761
rect 403 18659 437 18693
rect 403 18591 437 18625
rect 403 18523 437 18557
rect 403 18455 437 18489
rect 403 18387 437 18421
rect 403 18319 437 18353
rect 403 18251 437 18285
rect 403 18183 437 18217
rect 403 18115 437 18149
rect 403 18047 437 18081
rect 403 17979 437 18013
rect 403 17911 437 17945
rect 403 17843 437 17877
rect 403 17775 437 17809
rect 403 17707 437 17741
rect 403 17639 437 17673
rect 403 17571 437 17605
rect 403 17503 437 17537
rect 403 17435 437 17469
rect 403 17367 437 17401
rect 403 17299 437 17333
rect 403 17231 437 17265
rect 403 17163 437 17197
rect 403 17095 437 17129
rect 403 17027 437 17061
rect 403 16959 437 16993
rect 403 16891 437 16925
rect 403 16823 437 16857
rect 403 16755 437 16789
rect 403 16687 437 16721
rect 403 16619 437 16653
rect 403 16551 437 16585
rect 403 16483 437 16517
rect 403 16415 437 16449
rect 403 16347 437 16381
rect 403 16279 437 16313
rect 403 16211 437 16245
rect 403 16143 437 16177
rect 403 16075 437 16109
rect 403 16007 437 16041
rect 403 15939 437 15973
rect 403 15871 437 15905
rect 403 15803 437 15837
rect 403 15735 437 15769
rect 403 15667 437 15701
rect 403 15599 437 15633
rect 403 15531 437 15565
rect 403 15463 437 15497
rect 403 15395 437 15429
rect 403 15327 437 15361
rect 403 15259 437 15293
rect 403 15197 437 15225
rect 12423 21325 12457 21359
rect 12423 21257 12457 21291
rect 12423 21189 12457 21223
rect 12423 21121 12457 21155
rect 12423 21053 12457 21087
rect 12423 20985 12457 21019
rect 12423 20917 12457 20951
rect 12423 20849 12457 20883
rect 12423 20781 12457 20815
rect 12423 20713 12457 20747
rect 12423 20645 12457 20679
rect 12423 20577 12457 20611
rect 12423 20509 12457 20543
rect 12423 20441 12457 20475
rect 12423 20373 12457 20407
rect 12423 20305 12457 20339
rect 12423 20237 12457 20271
rect 12423 20169 12457 20203
rect 12423 20101 12457 20135
rect 12423 20033 12457 20067
rect 12423 19965 12457 19999
rect 12423 19897 12457 19931
rect 12423 19829 12457 19863
rect 12423 19761 12457 19795
rect 12423 19693 12457 19727
rect 12423 19625 12457 19659
rect 12423 19557 12457 19591
rect 12423 19489 12457 19523
rect 12423 19421 12457 19455
rect 12423 19353 12457 19387
rect 12423 19285 12457 19319
rect 12423 19217 12457 19251
rect 12423 19149 12457 19183
rect 12423 19081 12457 19115
rect 12423 19013 12457 19047
rect 12423 18945 12457 18979
rect 12423 18877 12457 18911
rect 12423 18809 12457 18843
rect 12423 18741 12457 18775
rect 12423 18673 12457 18707
rect 12423 18605 12457 18639
rect 12423 18537 12457 18571
rect 12423 18469 12457 18503
rect 12423 18401 12457 18435
rect 12423 18333 12457 18367
rect 12423 18265 12457 18299
rect 12423 18197 12457 18231
rect 12423 18129 12457 18163
rect 12423 18061 12457 18095
rect 12423 17993 12457 18027
rect 12423 17925 12457 17959
rect 12423 17857 12457 17891
rect 12423 17789 12457 17823
rect 12423 17721 12457 17755
rect 12423 17653 12457 17687
rect 12423 17585 12457 17619
rect 12423 17517 12457 17551
rect 12423 17449 12457 17483
rect 12423 17381 12457 17415
rect 12423 17313 12457 17347
rect 12423 17245 12457 17279
rect 12423 17177 12457 17211
rect 12423 17109 12457 17143
rect 12423 17041 12457 17075
rect 12423 16973 12457 17007
rect 12423 16905 12457 16939
rect 12423 16837 12457 16871
rect 12423 16769 12457 16803
rect 12423 16701 12457 16735
rect 12423 16633 12457 16667
rect 12423 16565 12457 16599
rect 12423 16497 12457 16531
rect 12423 16429 12457 16463
rect 12423 16361 12457 16395
rect 12423 16293 12457 16327
rect 12423 16225 12457 16259
rect 12423 16157 12457 16191
rect 12423 16089 12457 16123
rect 12423 16021 12457 16055
rect 12423 15953 12457 15987
rect 12423 15885 12457 15919
rect 12423 15817 12457 15851
rect 12423 15749 12457 15783
rect 12423 15681 12457 15715
rect 12423 15613 12457 15647
rect 12423 15545 12457 15579
rect 12423 15477 12457 15511
rect 12423 15409 12457 15443
rect 12423 15341 12457 15375
rect 12423 15273 12457 15307
rect 12423 15197 12457 15239
rect 403 15163 463 15197
rect 497 15163 531 15197
rect 565 15163 599 15197
rect 633 15163 667 15197
rect 701 15163 735 15197
rect 769 15163 803 15197
rect 837 15163 871 15197
rect 905 15163 939 15197
rect 973 15163 1007 15197
rect 1041 15163 1075 15197
rect 1109 15163 1143 15197
rect 1177 15163 1211 15197
rect 1245 15163 1279 15197
rect 1313 15163 1347 15197
rect 1381 15163 1415 15197
rect 1449 15163 1483 15197
rect 1517 15163 1551 15197
rect 1585 15163 1619 15197
rect 1653 15163 1687 15197
rect 1721 15163 1755 15197
rect 1789 15163 1823 15197
rect 1857 15163 1891 15197
rect 1925 15163 1959 15197
rect 1993 15163 2027 15197
rect 2061 15163 2095 15197
rect 2129 15163 2163 15197
rect 2197 15163 2231 15197
rect 2265 15163 2299 15197
rect 2333 15163 2367 15197
rect 2401 15163 2435 15197
rect 2469 15163 2503 15197
rect 2537 15163 2571 15197
rect 2605 15163 2639 15197
rect 2673 15163 2707 15197
rect 2741 15163 2775 15197
rect 2809 15163 2843 15197
rect 2877 15163 2911 15197
rect 2945 15163 2979 15197
rect 3013 15163 3047 15197
rect 3081 15163 3115 15197
rect 3149 15163 3183 15197
rect 3217 15163 3251 15197
rect 3285 15163 3319 15197
rect 3353 15163 3387 15197
rect 3421 15163 3455 15197
rect 3489 15163 3523 15197
rect 3557 15163 3591 15197
rect 3625 15163 3659 15197
rect 3693 15163 3727 15197
rect 3761 15163 3795 15197
rect 3829 15163 3863 15197
rect 3897 15163 3931 15197
rect 3965 15163 3999 15197
rect 4033 15163 4067 15197
rect 4101 15163 4135 15197
rect 4169 15163 4203 15197
rect 4237 15163 4271 15197
rect 4305 15163 4339 15197
rect 4373 15163 4407 15197
rect 4441 15163 4475 15197
rect 4509 15163 4543 15197
rect 4577 15163 4611 15197
rect 4645 15163 4679 15197
rect 4713 15163 4747 15197
rect 4781 15163 4815 15197
rect 4849 15163 4883 15197
rect 4917 15163 4951 15197
rect 4985 15163 5019 15197
rect 5053 15163 5087 15197
rect 5121 15163 5155 15197
rect 5189 15163 5223 15197
rect 5257 15163 5291 15197
rect 5325 15163 5359 15197
rect 5393 15163 5427 15197
rect 5461 15163 5495 15197
rect 5529 15163 5563 15197
rect 5597 15163 5631 15197
rect 5665 15163 5699 15197
rect 5733 15163 5767 15197
rect 5801 15163 5835 15197
rect 5869 15163 5903 15197
rect 5937 15163 5971 15197
rect 6005 15163 6039 15197
rect 6073 15163 6107 15197
rect 6141 15163 6175 15197
rect 6209 15163 6243 15197
rect 6277 15163 6311 15197
rect 6345 15163 6379 15197
rect 6413 15163 6447 15197
rect 6481 15163 6515 15197
rect 6549 15163 6583 15197
rect 6617 15163 6651 15197
rect 6685 15163 6719 15197
rect 6753 15163 6787 15197
rect 6821 15163 6855 15197
rect 6889 15163 6923 15197
rect 6957 15163 6991 15197
rect 7025 15163 7059 15197
rect 7093 15163 7127 15197
rect 7161 15163 7195 15197
rect 7229 15163 7263 15197
rect 7297 15163 7331 15197
rect 7365 15163 7399 15197
rect 7433 15163 7467 15197
rect 7501 15163 7535 15197
rect 7569 15163 7603 15197
rect 7637 15163 7671 15197
rect 7705 15163 7739 15197
rect 7773 15163 7807 15197
rect 7841 15163 7875 15197
rect 7909 15163 7943 15197
rect 7977 15163 8011 15197
rect 8045 15163 8079 15197
rect 8113 15163 8147 15197
rect 8181 15163 8215 15197
rect 8249 15163 8283 15197
rect 8317 15163 8351 15197
rect 8385 15163 8419 15197
rect 8453 15163 8487 15197
rect 8521 15163 8555 15197
rect 8589 15163 8623 15197
rect 8657 15163 8691 15197
rect 8725 15163 8759 15197
rect 8793 15163 8827 15197
rect 8861 15163 8895 15197
rect 8929 15163 8963 15197
rect 8997 15163 9031 15197
rect 9065 15163 9099 15197
rect 9133 15163 9167 15197
rect 9201 15163 9235 15197
rect 9269 15163 9303 15197
rect 9337 15163 9371 15197
rect 9405 15163 9439 15197
rect 9473 15163 9507 15197
rect 9541 15163 9575 15197
rect 9609 15163 9643 15197
rect 9677 15163 9711 15197
rect 9745 15163 9779 15197
rect 9813 15163 9847 15197
rect 9881 15163 9915 15197
rect 9949 15163 9983 15197
rect 10017 15163 10051 15197
rect 10085 15163 10119 15197
rect 10153 15163 10187 15197
rect 10221 15163 10255 15197
rect 10289 15163 10323 15197
rect 10357 15163 10391 15197
rect 10425 15163 10459 15197
rect 10493 15163 10527 15197
rect 10561 15163 10595 15197
rect 10629 15163 10663 15197
rect 10697 15163 10731 15197
rect 10765 15163 10799 15197
rect 10833 15163 10867 15197
rect 10901 15163 10935 15197
rect 10969 15163 11003 15197
rect 11037 15163 11071 15197
rect 11105 15163 11139 15197
rect 11173 15163 11207 15197
rect 11241 15163 11275 15197
rect 11309 15163 11343 15197
rect 11377 15163 11411 15197
rect 11445 15163 11479 15197
rect 11513 15163 11547 15197
rect 11581 15163 11615 15197
rect 11649 15163 11683 15197
rect 11717 15163 11751 15197
rect 11785 15163 11819 15197
rect 11853 15163 11887 15197
rect 11921 15163 11955 15197
rect 11989 15163 12023 15197
rect 12057 15163 12091 15197
rect 12125 15163 12159 15197
rect 12193 15163 12227 15197
rect 12261 15163 12295 15197
rect 12329 15163 12363 15197
rect 12397 15163 12457 15197
<< psubdiffcont >>
rect 458 13183 492 13217
rect 526 13183 560 13217
rect 594 13183 628 13217
rect 662 13183 696 13217
rect 730 13183 764 13217
rect 798 13183 832 13217
rect 866 13183 900 13217
rect 934 13183 968 13217
rect 1002 13183 1036 13217
rect 1070 13183 1104 13217
rect 1138 13183 1172 13217
rect 1206 13183 1240 13217
rect 1274 13183 1308 13217
rect 1342 13183 1376 13217
rect 1410 13183 1444 13217
rect 1478 13183 1512 13217
rect 1546 13183 1580 13217
rect 1614 13183 1648 13217
rect 1682 13183 1716 13217
rect 1750 13183 1784 13217
rect 1818 13183 1852 13217
rect 1886 13183 1920 13217
rect 1954 13183 1988 13217
rect 2022 13183 2056 13217
rect 2090 13183 2124 13217
rect 2158 13183 2192 13217
rect 2226 13183 2260 13217
rect 2294 13183 2328 13217
rect 2362 13183 2396 13217
rect 2430 13183 2464 13217
rect 2498 13183 2532 13217
rect 2566 13183 2600 13217
rect 2634 13183 2668 13217
rect 2702 13183 2736 13217
rect 2770 13183 2804 13217
rect 2838 13183 2872 13217
rect 2906 13183 2940 13217
rect 2974 13183 3008 13217
rect 3042 13183 3076 13217
rect 3110 13183 3144 13217
rect 3178 13183 3212 13217
rect 3246 13183 3280 13217
rect 3314 13183 3348 13217
rect 3382 13183 3416 13217
rect 3450 13183 3484 13217
rect 3518 13183 3552 13217
rect 3586 13183 3620 13217
rect 3654 13183 3688 13217
rect 3722 13183 3756 13217
rect 3790 13183 3824 13217
rect 3858 13183 3892 13217
rect 3926 13183 3960 13217
rect 3994 13183 4028 13217
rect 4062 13183 4096 13217
rect 4130 13183 4164 13217
rect 4198 13183 4232 13217
rect 4266 13183 4300 13217
rect 4334 13183 4368 13217
rect 4402 13183 4436 13217
rect 4470 13183 4504 13217
rect 4538 13183 4572 13217
rect 4606 13183 4640 13217
rect 4674 13183 4708 13217
rect 4742 13183 4776 13217
rect 4810 13183 4844 13217
rect 4878 13183 4912 13217
rect 4946 13183 4980 13217
rect 5014 13183 5048 13217
rect 5082 13183 5116 13217
rect 5150 13183 5184 13217
rect 5218 13183 5252 13217
rect 5286 13183 5320 13217
rect 5354 13183 5388 13217
rect 5422 13183 5456 13217
rect 5490 13183 5524 13217
rect 5558 13183 5592 13217
rect 5626 13183 5660 13217
rect 5694 13183 5728 13217
rect 5762 13183 5796 13217
rect 5830 13183 5864 13217
rect 5898 13183 5932 13217
rect 5966 13183 6000 13217
rect 6034 13183 6068 13217
rect 6102 13183 6136 13217
rect 6170 13183 6204 13217
rect 6238 13183 6272 13217
rect 6306 13183 6340 13217
rect 6374 13183 6408 13217
rect 6442 13183 6476 13217
rect 6510 13183 6544 13217
rect 6578 13183 6612 13217
rect 6646 13183 6680 13217
rect 6714 13183 6748 13217
rect 6782 13183 6816 13217
rect 6850 13183 6884 13217
rect 6918 13183 6952 13217
rect 6986 13183 7020 13217
rect 7054 13183 7088 13217
rect 7122 13183 7156 13217
rect 7190 13183 7224 13217
rect 7258 13183 7292 13217
rect 7326 13183 7360 13217
rect 7394 13183 7428 13217
rect 7462 13183 7496 13217
rect 7530 13183 7564 13217
rect 7598 13183 7632 13217
rect 7666 13183 7700 13217
rect 7734 13183 7768 13217
rect 7802 13183 7836 13217
rect 7870 13183 7904 13217
rect 7938 13183 7972 13217
rect 8006 13183 8040 13217
rect 8074 13183 8108 13217
rect 8142 13183 8176 13217
rect 8210 13183 8244 13217
rect 8278 13183 8312 13217
rect 8346 13183 8380 13217
rect 8414 13183 8448 13217
rect 8482 13183 8516 13217
rect 8550 13183 8584 13217
rect 8618 13183 8652 13217
rect 8686 13183 8720 13217
rect 8754 13183 8788 13217
rect 8822 13183 8856 13217
rect 8890 13183 8924 13217
rect 8958 13183 8992 13217
rect 9026 13183 9060 13217
rect 9094 13183 9128 13217
rect 9162 13183 9196 13217
rect 9230 13183 9264 13217
rect 9384 13183 9418 13217
rect 9452 13183 9486 13217
rect 9520 13183 9554 13217
rect 9588 13183 9622 13217
rect 9656 13183 9690 13217
rect 9724 13183 9758 13217
rect 9792 13183 9826 13217
rect 9860 13183 9894 13217
rect 9928 13183 9962 13217
rect 9996 13183 10030 13217
rect 10064 13183 10098 13217
rect 10132 13183 10166 13217
rect 10200 13183 10234 13217
rect 10268 13183 10302 13217
rect 10336 13183 10370 13217
rect 10404 13183 10438 13217
rect 10472 13183 10506 13217
rect 10540 13183 10574 13217
rect 10608 13183 10642 13217
rect 10676 13183 10710 13217
rect 10744 13183 10778 13217
rect 10812 13183 10846 13217
rect 10880 13183 10914 13217
rect 10948 13183 10982 13217
rect 11016 13183 11050 13217
rect 11084 13183 11118 13217
rect 11152 13183 11186 13217
rect 11220 13183 11254 13217
rect 11288 13183 11322 13217
rect 11356 13183 11390 13217
rect 11424 13183 11458 13217
rect 11492 13183 11526 13217
rect 383 13101 417 13135
rect 383 13033 417 13067
rect 383 12965 417 12999
rect 383 12897 417 12931
rect 383 12829 417 12863
rect 383 12761 417 12795
rect 383 12693 417 12727
rect 383 12625 417 12659
rect 383 12557 417 12591
rect 383 12489 417 12523
rect 383 12421 417 12455
rect 11573 13103 11607 13137
rect 11573 13035 11607 13069
rect 11573 12967 11607 13001
rect 11573 12899 11607 12933
rect 11573 12831 11607 12865
rect 11573 12763 11607 12797
rect 11573 12695 11607 12729
rect 11573 12627 11607 12661
rect 11573 12559 11607 12593
rect 11573 12491 11607 12525
rect 11573 12423 11607 12457
rect 383 12353 417 12387
rect 383 12285 417 12319
rect 2723 12313 2757 12347
rect 2903 12313 2937 12347
rect 5623 12303 5657 12337
rect 383 12217 417 12251
rect 5803 12303 5837 12337
rect 11573 12355 11607 12389
rect 11573 12287 11607 12321
rect 383 12149 417 12183
rect 383 12081 417 12115
rect 383 12013 417 12047
rect 383 11945 417 11979
rect 383 11877 417 11911
rect 383 11809 417 11843
rect 383 11741 417 11775
rect 383 11673 417 11707
rect 383 11605 417 11639
rect 383 11537 417 11571
rect 383 11469 417 11503
rect 383 11401 417 11435
rect 383 11333 417 11367
rect 383 11265 417 11299
rect 383 11197 417 11231
rect 383 11129 417 11163
rect 383 11061 417 11095
rect 383 10993 417 11027
rect 11573 12219 11607 12253
rect 11573 12151 11607 12185
rect 11573 12083 11607 12117
rect 11573 12015 11607 12049
rect 11573 11947 11607 11981
rect 11573 11879 11607 11913
rect 11573 11811 11607 11845
rect 11573 11743 11607 11777
rect 11573 11675 11607 11709
rect 11573 11607 11607 11641
rect 11573 11539 11607 11573
rect 11573 11471 11607 11505
rect 11573 11403 11607 11437
rect 11573 11335 11607 11369
rect 11573 11267 11607 11301
rect 11573 11199 11607 11233
rect 11573 11131 11607 11165
rect 11573 11063 11607 11097
rect 11644 10983 11678 11017
rect 11712 10983 11746 11017
rect 11780 10983 11814 11017
rect 11848 10983 11882 11017
rect 11916 10983 11950 11017
rect 11984 10983 12018 11017
rect 12052 10983 12086 11017
rect 12120 10983 12154 11017
rect 12188 10983 12222 11017
rect 12256 10983 12290 11017
rect 12324 10983 12358 11017
rect 12392 10983 12426 11017
rect 12460 10983 12494 11017
rect 12528 10983 12562 11017
rect 12596 10983 12630 11017
rect 12664 10983 12698 11017
rect 12732 10983 12766 11017
rect 12800 10983 12834 11017
rect 12868 10983 12902 11017
rect 12936 10983 12970 11017
rect 13004 10983 13038 11017
rect 13072 10983 13106 11017
rect 13140 10983 13174 11017
rect 13208 10983 13242 11017
rect 13276 10983 13310 11017
rect 13344 10983 13378 11017
rect 13412 10983 13446 11017
rect 13480 10983 13514 11017
rect 13548 10983 13582 11017
rect 13616 10983 13650 11017
rect 13684 10983 13718 11017
rect 13752 10983 13786 11017
rect 13820 10983 13854 11017
rect 13888 10983 13922 11017
rect 13956 10983 13990 11017
rect 14024 10983 14058 11017
rect 14092 10983 14126 11017
rect 14160 10983 14194 11017
rect 14228 10983 14262 11017
rect 14296 10983 14330 11017
rect 14364 10983 14398 11017
rect 14432 10983 14466 11017
rect 14500 10983 14534 11017
rect 14568 10983 14602 11017
rect 14636 10983 14670 11017
rect 14704 10983 14738 11017
rect 14772 10983 14806 11017
rect 14840 10983 14874 11017
rect 14908 10983 14942 11017
rect 14976 10983 15010 11017
rect 15044 10983 15078 11017
rect 15112 10983 15146 11017
rect 15180 10983 15214 11017
rect 15248 10983 15282 11017
rect 15316 10983 15350 11017
rect 15384 10983 15418 11017
rect 15452 10983 15486 11017
rect 15520 10983 15554 11017
rect 15588 10983 15622 11017
rect 15656 10983 15690 11017
rect 15724 10983 15758 11017
rect 15792 10983 15826 11017
rect 15860 10983 15894 11017
rect 15928 10983 15962 11017
rect 15996 10983 16030 11017
rect 16064 10983 16098 11017
rect 16132 10983 16166 11017
rect 16200 10983 16234 11017
rect 16268 10983 16302 11017
rect 16336 10983 16370 11017
rect 16404 10983 16438 11017
rect 16472 10983 16506 11017
rect 16540 10983 16574 11017
rect 16608 10983 16642 11017
rect 16676 10983 16710 11017
rect 16744 10983 16778 11017
rect 16812 10983 16846 11017
rect 16880 10983 16914 11017
rect 16948 10983 16982 11017
rect 17016 10983 17050 11017
rect 17084 10983 17118 11017
rect 17152 10983 17186 11017
rect 17220 10983 17254 11017
rect 17288 10983 17322 11017
rect 17356 10983 17390 11017
rect 17424 10983 17458 11017
rect 17492 10983 17526 11017
rect 17560 10983 17594 11017
rect 17628 10983 17662 11017
rect 17696 10983 17730 11017
rect 17764 10983 17798 11017
rect 17832 10983 17866 11017
rect 17900 10983 17934 11017
rect 17968 10983 18002 11017
rect 18036 10983 18070 11017
rect 18104 10983 18138 11017
rect 18172 10983 18206 11017
rect 18240 10983 18274 11017
rect 18308 10983 18342 11017
rect 18376 10983 18410 11017
rect 18444 10983 18478 11017
rect 18512 10983 18546 11017
rect 18580 10983 18614 11017
rect 18648 10983 18682 11017
rect 18716 10983 18750 11017
rect 18784 10983 18818 11017
rect 18852 10983 18886 11017
rect 18920 10983 18954 11017
rect 18988 10983 19022 11017
rect 19056 10983 19090 11017
rect 19124 10983 19158 11017
rect 19192 10983 19226 11017
rect 19260 10983 19294 11017
rect 19328 10983 19362 11017
rect 19396 10983 19430 11017
rect 19464 10983 19498 11017
rect 19532 10983 19566 11017
rect 19600 10983 19634 11017
rect 19668 10983 19702 11017
rect 19736 10983 19770 11017
rect 19804 10983 19838 11017
rect 19872 10983 19906 11017
rect 19940 10983 19974 11017
rect 20008 10983 20042 11017
rect 20076 10983 20110 11017
rect 20144 10983 20178 11017
rect 20212 10983 20246 11017
rect 20280 10983 20314 11017
rect 20348 10983 20382 11017
rect 20416 10983 20450 11017
rect 20484 10983 20518 11017
rect 20552 10983 20586 11017
rect 20620 10983 20654 11017
rect 20688 10983 20722 11017
rect 20756 10983 20790 11017
rect 20824 10983 20858 11017
rect 20892 10983 20926 11017
rect 20960 10983 20994 11017
rect 21028 10983 21062 11017
rect 21096 10983 21130 11017
rect 21164 10983 21198 11017
rect 21232 10983 21266 11017
rect 21300 10983 21334 11017
rect 21368 10983 21402 11017
rect 21436 10983 21470 11017
rect 21504 10983 21538 11017
rect 21572 10983 21606 11017
rect 21640 10983 21674 11017
rect 21708 10983 21742 11017
rect 21776 10983 21810 11017
rect 21844 10983 21878 11017
rect 21912 10983 21946 11017
rect 21980 10983 22014 11017
rect 22048 10983 22082 11017
rect 22116 10983 22150 11017
rect 22184 10983 22218 11017
rect 22252 10983 22286 11017
rect 22320 10983 22354 11017
rect 22388 10983 22422 11017
rect 383 10925 417 10959
rect 383 10857 417 10891
rect 383 10789 417 10823
rect 383 10721 417 10755
rect 383 10653 417 10687
rect 383 10585 417 10619
rect 383 10517 417 10551
rect 383 10449 417 10483
rect 22463 10913 22497 10947
rect 22463 10845 22497 10879
rect 22463 10777 22497 10811
rect 22463 10709 22497 10743
rect 22463 10641 22497 10675
rect 22463 10573 22497 10607
rect 22463 10505 22497 10539
rect 383 10381 417 10415
rect 383 10313 417 10347
rect 14323 10373 14357 10407
rect 22463 10437 22497 10471
rect 22463 10369 22497 10403
rect 383 10245 417 10279
rect 383 10177 417 10211
rect 383 10109 417 10143
rect 383 10041 417 10075
rect 383 9973 417 10007
rect 383 9905 417 9939
rect 383 9837 417 9871
rect 383 9769 417 9803
rect 383 9701 417 9735
rect 383 9633 417 9667
rect 383 9565 417 9599
rect 383 9497 417 9531
rect 383 9429 417 9463
rect 383 9361 417 9395
rect 383 9293 417 9327
rect 383 9225 417 9259
rect 383 9157 417 9191
rect 383 9089 417 9123
rect 383 9021 417 9055
rect 383 8953 417 8987
rect 383 8885 417 8919
rect 383 8817 417 8851
rect 383 8749 417 8783
rect 383 8681 417 8715
rect 383 8613 417 8647
rect 383 8545 417 8579
rect 383 8477 417 8511
rect 383 8409 417 8443
rect 383 8341 417 8375
rect 383 8273 417 8307
rect 383 8205 417 8239
rect 383 8137 417 8171
rect 383 8069 417 8103
rect 383 8001 417 8035
rect 383 7933 417 7967
rect 383 7865 417 7899
rect 383 7797 417 7831
rect 383 7729 417 7763
rect 383 7661 417 7695
rect 383 7593 417 7627
rect 383 7525 417 7559
rect 383 7457 417 7491
rect 383 7389 417 7423
rect 383 7321 417 7355
rect 383 7253 417 7287
rect 383 7185 417 7219
rect 383 7117 417 7151
rect 383 7049 417 7083
rect 383 6981 417 7015
rect 383 6913 417 6947
rect 383 6845 417 6879
rect 383 6777 417 6811
rect 383 6709 417 6743
rect 383 6641 417 6675
rect 383 6573 417 6607
rect 383 6505 417 6539
rect 383 6437 417 6471
rect 383 6369 417 6403
rect 383 6301 417 6335
rect 383 6233 417 6267
rect 383 6165 417 6199
rect 383 6097 417 6131
rect 383 6029 417 6063
rect 383 5961 417 5995
rect 22463 10301 22497 10335
rect 22463 10233 22497 10267
rect 22463 10165 22497 10199
rect 22463 10097 22497 10131
rect 22463 10029 22497 10063
rect 22463 9961 22497 9995
rect 22463 9893 22497 9927
rect 22463 9825 22497 9859
rect 22463 9757 22497 9791
rect 22463 9689 22497 9723
rect 22463 9621 22497 9655
rect 22463 9553 22497 9587
rect 22463 9485 22497 9519
rect 22463 9417 22497 9451
rect 22463 9349 22497 9383
rect 22463 9281 22497 9315
rect 22463 9213 22497 9247
rect 22463 9145 22497 9179
rect 22463 9077 22497 9111
rect 22463 9009 22497 9043
rect 22463 8941 22497 8975
rect 22463 8873 22497 8907
rect 22463 8805 22497 8839
rect 22463 8737 22497 8771
rect 22463 8669 22497 8703
rect 22463 8601 22497 8635
rect 22463 8533 22497 8567
rect 22463 8465 22497 8499
rect 22463 8397 22497 8431
rect 22463 8329 22497 8363
rect 22463 8261 22497 8295
rect 22463 8193 22497 8227
rect 22463 8125 22497 8159
rect 22463 8057 22497 8091
rect 22463 7989 22497 8023
rect 22463 7921 22497 7955
rect 22463 7853 22497 7887
rect 22463 7785 22497 7819
rect 22463 7717 22497 7751
rect 22463 7649 22497 7683
rect 22463 7581 22497 7615
rect 22463 7513 22497 7547
rect 22463 7445 22497 7479
rect 22463 7377 22497 7411
rect 22463 7309 22497 7343
rect 22463 7241 22497 7275
rect 22463 7173 22497 7207
rect 22463 7105 22497 7139
rect 22463 7037 22497 7071
rect 22463 6969 22497 7003
rect 22463 6901 22497 6935
rect 22463 6833 22497 6867
rect 22463 6765 22497 6799
rect 22463 6697 22497 6731
rect 22463 6629 22497 6663
rect 22463 6561 22497 6595
rect 22463 6493 22497 6527
rect 22463 6425 22497 6459
rect 22463 6357 22497 6391
rect 22463 6289 22497 6323
rect 22463 6221 22497 6255
rect 22463 6153 22497 6187
rect 22463 6085 22497 6119
rect 22463 6017 22497 6051
rect 22463 5949 22497 5983
rect 383 5893 417 5927
rect 383 5825 417 5859
rect 383 5757 417 5791
rect 1623 5843 1657 5877
rect 22463 5881 22497 5915
rect 22463 5813 22497 5847
rect 383 5689 417 5723
rect 383 5621 417 5655
rect 383 5553 417 5587
rect 383 5485 417 5519
rect 383 5417 417 5451
rect 383 5349 417 5383
rect 383 5281 417 5315
rect 383 5213 417 5247
rect 383 5145 417 5179
rect 383 5077 417 5111
rect 383 5009 417 5043
rect 383 4941 417 4975
rect 383 4873 417 4907
rect 383 4805 417 4839
rect 383 4737 417 4771
rect 383 4669 417 4703
rect 383 4601 417 4635
rect 383 4533 417 4567
rect 383 4465 417 4499
rect 383 4397 417 4431
rect 383 4329 417 4363
rect 383 4261 417 4295
rect 383 4193 417 4227
rect 383 4125 417 4159
rect 383 4057 417 4091
rect 383 3989 417 4023
rect 383 3921 417 3955
rect 383 3853 417 3887
rect 383 3785 417 3819
rect 383 3717 417 3751
rect 383 3649 417 3683
rect 383 3581 417 3615
rect 383 3513 417 3547
rect 383 3445 417 3479
rect 383 3377 417 3411
rect 383 3309 417 3343
rect 383 3241 417 3275
rect 383 3173 417 3207
rect 383 3105 417 3139
rect 383 3037 417 3071
rect 383 2969 417 3003
rect 383 2901 417 2935
rect 383 2833 417 2867
rect 383 2765 417 2799
rect 383 2697 417 2731
rect 383 2629 417 2663
rect 383 2561 417 2595
rect 383 2493 417 2527
rect 383 2425 417 2459
rect 383 2357 417 2391
rect 383 2289 417 2323
rect 383 2221 417 2255
rect 383 2153 417 2187
rect 383 2085 417 2119
rect 383 2017 417 2051
rect 383 1949 417 1983
rect 383 1881 417 1915
rect 383 1813 417 1847
rect 383 1745 417 1779
rect 383 1677 417 1711
rect 383 1609 417 1643
rect 383 1541 417 1575
rect 383 1473 417 1507
rect 383 1405 417 1439
rect 383 1337 417 1371
rect 383 1269 417 1303
rect 383 1201 417 1235
rect 383 1133 417 1167
rect 383 1065 417 1099
rect 383 997 417 1031
rect 383 929 417 963
rect 383 861 417 895
rect 383 793 417 827
rect 383 725 417 759
rect 383 657 417 691
rect 383 589 417 623
rect 383 521 417 555
rect 383 453 417 487
rect 383 385 417 419
rect 383 317 417 351
rect 383 249 417 283
rect 383 181 417 215
rect 383 113 417 147
rect 383 45 417 79
rect 383 -23 417 11
rect 383 -91 417 -57
rect 383 -159 417 -125
rect 383 -227 417 -193
rect 383 -295 417 -261
rect 383 -363 417 -329
rect 22463 5745 22497 5779
rect 22463 5677 22497 5711
rect 22463 5609 22497 5643
rect 22463 5541 22497 5575
rect 22463 5473 22497 5507
rect 22463 5405 22497 5439
rect 22463 5337 22497 5371
rect 22463 5269 22497 5303
rect 22463 5201 22497 5235
rect 22463 5133 22497 5167
rect 22463 5065 22497 5099
rect 22463 4997 22497 5031
rect 22463 4929 22497 4963
rect 22463 4861 22497 4895
rect 22463 4793 22497 4827
rect 22463 4725 22497 4759
rect 22463 4657 22497 4691
rect 22463 4589 22497 4623
rect 22463 4521 22497 4555
rect 22463 4453 22497 4487
rect 22463 4385 22497 4419
rect 22463 4317 22497 4351
rect 22463 4249 22497 4283
rect 22463 4181 22497 4215
rect 22463 4113 22497 4147
rect 22463 4045 22497 4079
rect 22463 3977 22497 4011
rect 22463 3909 22497 3943
rect 22463 3841 22497 3875
rect 22463 3773 22497 3807
rect 22463 3705 22497 3739
rect 22463 3637 22497 3671
rect 22463 3569 22497 3603
rect 22463 3501 22497 3535
rect 22463 3433 22497 3467
rect 22463 3365 22497 3399
rect 22463 3297 22497 3331
rect 22463 3229 22497 3263
rect 22463 3161 22497 3195
rect 22463 3093 22497 3127
rect 22463 3025 22497 3059
rect 22463 2957 22497 2991
rect 22463 2889 22497 2923
rect 22463 2821 22497 2855
rect 22463 2753 22497 2787
rect 22463 2685 22497 2719
rect 22463 2617 22497 2651
rect 22463 2549 22497 2583
rect 22463 2481 22497 2515
rect 22463 2413 22497 2447
rect 22463 2345 22497 2379
rect 22463 2277 22497 2311
rect 22463 2209 22497 2243
rect 22463 2141 22497 2175
rect 22463 2073 22497 2107
rect 22463 2005 22497 2039
rect 22463 1937 22497 1971
rect 22463 1869 22497 1903
rect 22463 1801 22497 1835
rect 22463 1733 22497 1767
rect 22463 1665 22497 1699
rect 22463 1597 22497 1631
rect 22463 1529 22497 1563
rect 22463 1461 22497 1495
rect 22463 1393 22497 1427
rect 22463 1325 22497 1359
rect 22463 1257 22497 1291
rect 22463 1189 22497 1223
rect 22463 1121 22497 1155
rect 22463 1053 22497 1087
rect 22463 985 22497 1019
rect 22463 917 22497 951
rect 22463 849 22497 883
rect 22463 781 22497 815
rect 22463 713 22497 747
rect 22463 645 22497 679
rect 22463 577 22497 611
rect 22463 509 22497 543
rect 22463 441 22497 475
rect 22463 373 22497 407
rect 22463 305 22497 339
rect 22463 237 22497 271
rect 22463 169 22497 203
rect 22463 101 22497 135
rect 22463 33 22497 67
rect 22463 -35 22497 -1
rect 22463 -103 22497 -69
rect 22463 -171 22497 -137
rect 22463 -239 22497 -205
rect 22463 -307 22497 -273
rect 383 -431 417 -397
rect 22463 -375 22497 -341
rect 383 -499 417 -465
rect 383 -567 417 -533
rect 1533 -527 1567 -493
rect 1713 -527 1747 -493
rect 19173 -457 19207 -423
rect 21143 -467 21177 -433
rect 21513 -467 21547 -433
rect 22463 -443 22497 -409
rect 22463 -511 22497 -477
rect 22463 -579 22497 -545
rect 383 -635 417 -601
rect 22463 -647 22497 -613
rect 475 -717 509 -683
rect 543 -717 577 -683
rect 611 -717 645 -683
rect 679 -717 713 -683
rect 747 -717 781 -683
rect 815 -717 849 -683
rect 883 -717 917 -683
rect 951 -717 985 -683
rect 1019 -717 1053 -683
rect 1087 -717 1121 -683
rect 1155 -717 1189 -683
rect 1223 -717 1257 -683
rect 1291 -717 1325 -683
rect 1359 -717 1393 -683
rect 1427 -717 1461 -683
rect 1495 -717 1529 -683
rect 1563 -717 1597 -683
rect 1631 -717 1665 -683
rect 1699 -717 1733 -683
rect 1767 -717 1801 -683
rect 1835 -717 1869 -683
rect 1903 -717 1937 -683
rect 1971 -717 2005 -683
rect 2039 -717 2073 -683
rect 2107 -717 2141 -683
rect 2175 -717 2209 -683
rect 2243 -717 2277 -683
rect 2311 -717 2345 -683
rect 2379 -717 2413 -683
rect 2447 -717 2481 -683
rect 2515 -717 2549 -683
rect 2583 -717 2617 -683
rect 2651 -717 2685 -683
rect 2719 -717 2753 -683
rect 2787 -717 2821 -683
rect 2855 -717 2889 -683
rect 2923 -717 2957 -683
rect 2991 -717 3025 -683
rect 3059 -717 3093 -683
rect 3127 -717 3161 -683
rect 3195 -717 3229 -683
rect 3263 -717 3297 -683
rect 3331 -717 3365 -683
rect 3399 -717 3433 -683
rect 3467 -717 3501 -683
rect 3535 -717 3569 -683
rect 3603 -717 3637 -683
rect 3671 -717 3705 -683
rect 3739 -717 3773 -683
rect 3807 -717 3841 -683
rect 3875 -717 3909 -683
rect 3943 -717 3977 -683
rect 4011 -717 4045 -683
rect 4079 -717 4113 -683
rect 4147 -717 4181 -683
rect 4215 -717 4249 -683
rect 4283 -717 4317 -683
rect 4351 -717 4385 -683
rect 4419 -717 4453 -683
rect 4487 -717 4521 -683
rect 4555 -717 4589 -683
rect 4623 -717 4657 -683
rect 4691 -717 4725 -683
rect 4759 -717 4793 -683
rect 4827 -717 4861 -683
rect 4895 -717 4929 -683
rect 4963 -717 4997 -683
rect 5031 -717 5065 -683
rect 5099 -717 5133 -683
rect 5167 -717 5201 -683
rect 5235 -717 5269 -683
rect 5303 -717 5337 -683
rect 5371 -717 5405 -683
rect 5439 -717 5473 -683
rect 5507 -717 5541 -683
rect 5575 -717 5609 -683
rect 5643 -717 5677 -683
rect 5711 -717 5745 -683
rect 5779 -717 5813 -683
rect 5847 -717 5881 -683
rect 5915 -717 5949 -683
rect 5983 -717 6017 -683
rect 6051 -717 6085 -683
rect 6119 -717 6153 -683
rect 6187 -717 6221 -683
rect 6255 -717 6289 -683
rect 6323 -717 6357 -683
rect 6391 -717 6425 -683
rect 6459 -717 6493 -683
rect 6527 -717 6561 -683
rect 6595 -717 6629 -683
rect 6663 -717 6697 -683
rect 6731 -717 6765 -683
rect 6799 -717 6833 -683
rect 6867 -717 6901 -683
rect 6935 -717 6969 -683
rect 7003 -717 7037 -683
rect 7071 -717 7105 -683
rect 7139 -717 7173 -683
rect 7207 -717 7241 -683
rect 7275 -717 7309 -683
rect 7343 -717 7377 -683
rect 7411 -717 7445 -683
rect 7479 -717 7513 -683
rect 7547 -717 7581 -683
rect 7615 -717 7649 -683
rect 7683 -717 7717 -683
rect 7751 -717 7785 -683
rect 7819 -717 7853 -683
rect 7887 -717 7921 -683
rect 7955 -717 7989 -683
rect 8023 -717 8057 -683
rect 8091 -717 8125 -683
rect 8159 -717 8193 -683
rect 8227 -717 8261 -683
rect 8295 -717 8329 -683
rect 8363 -717 8397 -683
rect 8431 -717 8465 -683
rect 8499 -717 8533 -683
rect 8567 -717 8601 -683
rect 8635 -717 8669 -683
rect 8703 -717 8737 -683
rect 8771 -717 8805 -683
rect 8839 -717 8873 -683
rect 8907 -717 8941 -683
rect 8975 -717 9009 -683
rect 9043 -717 9077 -683
rect 9111 -717 9145 -683
rect 9179 -717 9213 -683
rect 9247 -717 9281 -683
rect 9315 -717 9349 -683
rect 9383 -717 9417 -683
rect 9451 -717 9485 -683
rect 9519 -717 9553 -683
rect 9587 -717 9621 -683
rect 9655 -717 9689 -683
rect 9723 -717 9757 -683
rect 9791 -717 9825 -683
rect 9859 -717 9893 -683
rect 9927 -717 9961 -683
rect 9995 -717 10029 -683
rect 10063 -717 10097 -683
rect 10131 -717 10165 -683
rect 10199 -717 10233 -683
rect 10267 -717 10301 -683
rect 10335 -717 10369 -683
rect 10403 -717 10437 -683
rect 10471 -717 10505 -683
rect 10539 -717 10573 -683
rect 10607 -717 10641 -683
rect 10675 -717 10709 -683
rect 10743 -717 10777 -683
rect 10811 -717 10845 -683
rect 10879 -717 10913 -683
rect 10947 -717 10981 -683
rect 11015 -717 11049 -683
rect 11083 -717 11117 -683
rect 11151 -717 11185 -683
rect 11219 -717 11253 -683
rect 11287 -717 11321 -683
rect 11355 -717 11389 -683
rect 11423 -717 11457 -683
rect 11491 -717 11525 -683
rect 11559 -717 11593 -683
rect 11627 -717 11661 -683
rect 11695 -717 11729 -683
rect 11763 -717 11797 -683
rect 11831 -717 11865 -683
rect 11899 -717 11933 -683
rect 11967 -717 12001 -683
rect 12035 -717 12069 -683
rect 12103 -717 12137 -683
rect 12171 -717 12205 -683
rect 12239 -717 12273 -683
rect 12307 -717 12341 -683
rect 12375 -717 12409 -683
rect 12443 -717 12477 -683
rect 12511 -717 12545 -683
rect 12579 -717 12613 -683
rect 12647 -717 12681 -683
rect 12715 -717 12749 -683
rect 12783 -717 12817 -683
rect 12851 -717 12885 -683
rect 12919 -717 12953 -683
rect 12987 -717 13021 -683
rect 13055 -717 13089 -683
rect 13123 -717 13157 -683
rect 13191 -717 13225 -683
rect 13259 -717 13293 -683
rect 13327 -717 13361 -683
rect 13395 -717 13429 -683
rect 13463 -717 13497 -683
rect 13531 -717 13565 -683
rect 13599 -717 13633 -683
rect 13667 -717 13701 -683
rect 13735 -717 13769 -683
rect 13803 -717 13837 -683
rect 13871 -717 13905 -683
rect 13939 -717 13973 -683
rect 14007 -717 14041 -683
rect 14075 -717 14109 -683
rect 14143 -717 14177 -683
rect 14211 -717 14245 -683
rect 14279 -717 14313 -683
rect 14347 -717 14381 -683
rect 14415 -717 14449 -683
rect 14483 -717 14517 -683
rect 14551 -717 14585 -683
rect 14619 -717 14653 -683
rect 14687 -717 14721 -683
rect 14755 -717 14789 -683
rect 14823 -717 14857 -683
rect 14891 -717 14925 -683
rect 14959 -717 14993 -683
rect 15027 -717 15061 -683
rect 15095 -717 15129 -683
rect 15163 -717 15197 -683
rect 15231 -717 15265 -683
rect 15299 -717 15333 -683
rect 15367 -717 15401 -683
rect 15435 -717 15469 -683
rect 15503 -717 15537 -683
rect 15571 -717 15605 -683
rect 15639 -717 15673 -683
rect 15707 -717 15741 -683
rect 15775 -717 15809 -683
rect 15843 -717 15877 -683
rect 15911 -717 15945 -683
rect 15979 -717 16013 -683
rect 16047 -717 16081 -683
rect 16115 -717 16149 -683
rect 16183 -717 16217 -683
rect 16251 -717 16285 -683
rect 16319 -717 16353 -683
rect 16387 -717 16421 -683
rect 16455 -717 16489 -683
rect 16523 -717 16557 -683
rect 16591 -717 16625 -683
rect 16659 -717 16693 -683
rect 16727 -717 16761 -683
rect 16795 -717 16829 -683
rect 16863 -717 16897 -683
rect 16931 -717 16965 -683
rect 16999 -717 17033 -683
rect 17067 -717 17101 -683
rect 17135 -717 17169 -683
rect 17203 -717 17237 -683
rect 17271 -717 17305 -683
rect 17339 -717 17373 -683
rect 17407 -717 17441 -683
rect 17475 -717 17509 -683
rect 17543 -717 17577 -683
rect 17611 -717 17645 -683
rect 17679 -717 17713 -683
rect 17747 -717 17781 -683
rect 17815 -717 17849 -683
rect 17883 -717 17917 -683
rect 17951 -717 17985 -683
rect 18019 -717 18053 -683
rect 18087 -717 18121 -683
rect 18155 -717 18189 -683
rect 18223 -717 18257 -683
rect 18291 -717 18325 -683
rect 18359 -717 18393 -683
rect 18427 -717 18461 -683
rect 18495 -717 18529 -683
rect 18563 -717 18597 -683
rect 18631 -717 18665 -683
rect 18699 -717 18733 -683
rect 18767 -717 18801 -683
rect 18835 -717 18869 -683
rect 18903 -717 18937 -683
rect 18971 -717 19005 -683
rect 19039 -717 19073 -683
rect 19107 -717 19141 -683
rect 19175 -717 19209 -683
rect 19243 -717 19277 -683
rect 19311 -717 19345 -683
rect 19379 -717 19413 -683
rect 19447 -717 19481 -683
rect 19515 -717 19549 -683
rect 19583 -717 19617 -683
rect 19651 -717 19685 -683
rect 19719 -717 19753 -683
rect 19787 -717 19821 -683
rect 19855 -717 19889 -683
rect 19923 -717 19957 -683
rect 19991 -717 20025 -683
rect 20059 -717 20093 -683
rect 20127 -717 20161 -683
rect 20195 -717 20229 -683
rect 20263 -717 20297 -683
rect 20331 -717 20365 -683
rect 20399 -717 20433 -683
rect 20467 -717 20501 -683
rect 20535 -717 20569 -683
rect 20603 -717 20637 -683
rect 20671 -717 20705 -683
rect 20739 -717 20773 -683
rect 20807 -717 20841 -683
rect 20875 -717 20909 -683
rect 20943 -717 20977 -683
rect 21011 -717 21045 -683
rect 21079 -717 21113 -683
rect 21147 -717 21181 -683
rect 21215 -717 21249 -683
rect 21283 -717 21317 -683
rect 21351 -717 21385 -683
rect 21419 -717 21453 -683
rect 21487 -717 21521 -683
rect 21555 -717 21589 -683
rect 21623 -717 21657 -683
rect 21691 -717 21725 -683
rect 21759 -717 21793 -683
rect 21827 -717 21861 -683
rect 21895 -717 21929 -683
rect 21963 -717 21997 -683
rect 22031 -717 22065 -683
rect 22099 -717 22133 -683
rect 22167 -717 22201 -683
rect 22235 -717 22269 -683
rect 22303 -717 22337 -683
rect 22371 -717 22405 -683
<< nsubdiffcont >>
rect 403 21753 437 21787
rect 540 21783 574 21817
rect 608 21783 642 21817
rect 676 21783 710 21817
rect 744 21783 778 21817
rect 812 21783 846 21817
rect 880 21783 914 21817
rect 948 21783 982 21817
rect 1016 21783 1050 21817
rect 1084 21783 1118 21817
rect 1152 21783 1186 21817
rect 1220 21783 1254 21817
rect 1288 21783 1322 21817
rect 1356 21783 1390 21817
rect 1424 21783 1458 21817
rect 1492 21783 1526 21817
rect 1560 21783 1594 21817
rect 1628 21783 1662 21817
rect 1696 21783 1730 21817
rect 1764 21783 1798 21817
rect 1832 21783 1866 21817
rect 1900 21783 1934 21817
rect 1968 21783 2002 21817
rect 2036 21783 2070 21817
rect 2104 21783 2138 21817
rect 2172 21783 2206 21817
rect 2240 21783 2274 21817
rect 2308 21783 2342 21817
rect 2376 21783 2410 21817
rect 2444 21783 2478 21817
rect 2512 21783 2546 21817
rect 2580 21783 2614 21817
rect 2648 21783 2682 21817
rect 2716 21783 2750 21817
rect 2784 21783 2818 21817
rect 2852 21783 2886 21817
rect 2920 21783 2954 21817
rect 2988 21783 3022 21817
rect 3056 21783 3090 21817
rect 3124 21783 3158 21817
rect 3192 21783 3226 21817
rect 3260 21783 3294 21817
rect 3328 21783 3362 21817
rect 3396 21783 3430 21817
rect 3464 21783 3498 21817
rect 3532 21783 3566 21817
rect 3600 21783 3634 21817
rect 3668 21783 3702 21817
rect 3736 21783 3770 21817
rect 3804 21783 3838 21817
rect 3872 21783 3906 21817
rect 3940 21783 3974 21817
rect 4008 21783 4042 21817
rect 4076 21783 4110 21817
rect 4144 21783 4178 21817
rect 4212 21783 4246 21817
rect 4280 21783 4314 21817
rect 4348 21783 4382 21817
rect 4416 21783 4450 21817
rect 4484 21783 4518 21817
rect 4552 21783 4586 21817
rect 4620 21783 4654 21817
rect 4688 21783 4722 21817
rect 4756 21783 4790 21817
rect 4824 21783 4858 21817
rect 4892 21783 4926 21817
rect 4960 21783 4994 21817
rect 5028 21783 5062 21817
rect 5096 21783 5130 21817
rect 5164 21783 5198 21817
rect 5232 21783 5266 21817
rect 5300 21783 5334 21817
rect 5368 21783 5402 21817
rect 5436 21783 5470 21817
rect 5504 21783 5538 21817
rect 5572 21783 5606 21817
rect 5640 21783 5674 21817
rect 5708 21783 5742 21817
rect 5776 21783 5810 21817
rect 5844 21783 5878 21817
rect 5912 21783 5946 21817
rect 5980 21783 6014 21817
rect 6048 21783 6082 21817
rect 6116 21783 6150 21817
rect 6184 21783 6218 21817
rect 6252 21783 6286 21817
rect 6320 21783 6354 21817
rect 6388 21783 6422 21817
rect 6456 21783 6490 21817
rect 6524 21783 6558 21817
rect 6592 21783 6626 21817
rect 6660 21783 6694 21817
rect 6728 21783 6762 21817
rect 6796 21783 6830 21817
rect 6864 21783 6898 21817
rect 6932 21783 6966 21817
rect 7000 21783 7034 21817
rect 7068 21783 7102 21817
rect 7136 21783 7170 21817
rect 7204 21783 7238 21817
rect 7272 21783 7306 21817
rect 7340 21783 7374 21817
rect 7408 21783 7442 21817
rect 7476 21783 7510 21817
rect 7544 21783 7578 21817
rect 7612 21783 7646 21817
rect 7680 21783 7714 21817
rect 7748 21783 7782 21817
rect 7816 21783 7850 21817
rect 7884 21783 7918 21817
rect 7952 21783 7986 21817
rect 8020 21783 8054 21817
rect 8088 21783 8122 21817
rect 8156 21783 8190 21817
rect 8224 21783 8258 21817
rect 8292 21783 8326 21817
rect 8360 21783 8394 21817
rect 8428 21783 8462 21817
rect 8496 21783 8530 21817
rect 8564 21783 8598 21817
rect 8632 21783 8666 21817
rect 8700 21783 8734 21817
rect 8768 21783 8802 21817
rect 8836 21783 8870 21817
rect 8904 21783 8938 21817
rect 8972 21783 9006 21817
rect 9040 21783 9074 21817
rect 9108 21783 9142 21817
rect 9176 21783 9210 21817
rect 9244 21783 9278 21817
rect 9312 21783 9346 21817
rect 9380 21783 9414 21817
rect 9448 21783 9482 21817
rect 9516 21783 9550 21817
rect 9584 21783 9618 21817
rect 9652 21783 9686 21817
rect 9720 21783 9754 21817
rect 9788 21783 9822 21817
rect 9856 21783 9890 21817
rect 9924 21783 9958 21817
rect 9992 21783 10026 21817
rect 10060 21783 10094 21817
rect 10128 21783 10162 21817
rect 10196 21783 10230 21817
rect 10264 21783 10298 21817
rect 10332 21783 10366 21817
rect 10400 21783 10434 21817
rect 10468 21783 10502 21817
rect 10536 21783 10570 21817
rect 10604 21783 10638 21817
rect 10672 21783 10706 21817
rect 10740 21783 10774 21817
rect 10808 21783 10842 21817
rect 10876 21783 10910 21817
rect 10944 21783 10978 21817
rect 11012 21783 11046 21817
rect 11080 21783 11114 21817
rect 11148 21783 11182 21817
rect 11216 21783 11250 21817
rect 11284 21783 11318 21817
rect 11352 21783 11386 21817
rect 11420 21783 11454 21817
rect 11488 21783 11522 21817
rect 11556 21783 11590 21817
rect 11624 21783 11658 21817
rect 11692 21783 11726 21817
rect 11760 21783 11794 21817
rect 11828 21783 11862 21817
rect 11896 21783 11930 21817
rect 11964 21783 11998 21817
rect 12032 21783 12066 21817
rect 12100 21783 12134 21817
rect 12168 21783 12202 21817
rect 12236 21783 12270 21817
rect 12304 21783 12338 21817
rect 403 21685 437 21719
rect 403 21617 437 21651
rect 403 21549 437 21583
rect 403 21481 437 21515
rect 12423 21699 12457 21733
rect 12423 21631 12457 21665
rect 12423 21563 12457 21597
rect 12423 21495 12457 21529
rect 403 21413 437 21447
rect 1075 21408 1109 21442
rect 1143 21408 1177 21442
rect 1211 21408 1245 21442
rect 7055 21403 7089 21437
rect 7123 21403 7157 21437
rect 7191 21403 7225 21437
rect 403 21345 437 21379
rect 12423 21427 12457 21461
rect 403 21277 437 21311
rect 403 21209 437 21243
rect 403 21141 437 21175
rect 403 21073 437 21107
rect 403 21005 437 21039
rect 403 20937 437 20971
rect 403 20869 437 20903
rect 403 20801 437 20835
rect 403 20733 437 20767
rect 403 20665 437 20699
rect 403 20597 437 20631
rect 403 20529 437 20563
rect 403 20461 437 20495
rect 403 20393 437 20427
rect 403 20325 437 20359
rect 403 20257 437 20291
rect 403 20189 437 20223
rect 403 20121 437 20155
rect 403 20053 437 20087
rect 403 19985 437 20019
rect 403 19917 437 19951
rect 403 19849 437 19883
rect 403 19781 437 19815
rect 403 19713 437 19747
rect 403 19645 437 19679
rect 403 19577 437 19611
rect 403 19509 437 19543
rect 403 19441 437 19475
rect 403 19373 437 19407
rect 403 19305 437 19339
rect 403 19237 437 19271
rect 403 19169 437 19203
rect 403 19101 437 19135
rect 403 19033 437 19067
rect 403 18965 437 18999
rect 403 18897 437 18931
rect 403 18829 437 18863
rect 403 18761 437 18795
rect 403 18693 437 18727
rect 403 18625 437 18659
rect 403 18557 437 18591
rect 403 18489 437 18523
rect 403 18421 437 18455
rect 403 18353 437 18387
rect 403 18285 437 18319
rect 403 18217 437 18251
rect 403 18149 437 18183
rect 403 18081 437 18115
rect 403 18013 437 18047
rect 403 17945 437 17979
rect 403 17877 437 17911
rect 403 17809 437 17843
rect 403 17741 437 17775
rect 403 17673 437 17707
rect 403 17605 437 17639
rect 403 17537 437 17571
rect 403 17469 437 17503
rect 403 17401 437 17435
rect 403 17333 437 17367
rect 403 17265 437 17299
rect 403 17197 437 17231
rect 403 17129 437 17163
rect 403 17061 437 17095
rect 403 16993 437 17027
rect 403 16925 437 16959
rect 403 16857 437 16891
rect 403 16789 437 16823
rect 403 16721 437 16755
rect 403 16653 437 16687
rect 403 16585 437 16619
rect 403 16517 437 16551
rect 403 16449 437 16483
rect 403 16381 437 16415
rect 403 16313 437 16347
rect 403 16245 437 16279
rect 403 16177 437 16211
rect 403 16109 437 16143
rect 403 16041 437 16075
rect 403 15973 437 16007
rect 403 15905 437 15939
rect 403 15837 437 15871
rect 403 15769 437 15803
rect 403 15701 437 15735
rect 403 15633 437 15667
rect 403 15565 437 15599
rect 403 15497 437 15531
rect 403 15429 437 15463
rect 403 15361 437 15395
rect 403 15293 437 15327
rect 403 15225 437 15259
rect 12423 21359 12457 21393
rect 12423 21291 12457 21325
rect 12423 21223 12457 21257
rect 12423 21155 12457 21189
rect 12423 21087 12457 21121
rect 12423 21019 12457 21053
rect 12423 20951 12457 20985
rect 12423 20883 12457 20917
rect 12423 20815 12457 20849
rect 12423 20747 12457 20781
rect 12423 20679 12457 20713
rect 12423 20611 12457 20645
rect 12423 20543 12457 20577
rect 12423 20475 12457 20509
rect 12423 20407 12457 20441
rect 12423 20339 12457 20373
rect 12423 20271 12457 20305
rect 12423 20203 12457 20237
rect 12423 20135 12457 20169
rect 12423 20067 12457 20101
rect 12423 19999 12457 20033
rect 12423 19931 12457 19965
rect 12423 19863 12457 19897
rect 12423 19795 12457 19829
rect 12423 19727 12457 19761
rect 12423 19659 12457 19693
rect 12423 19591 12457 19625
rect 12423 19523 12457 19557
rect 12423 19455 12457 19489
rect 12423 19387 12457 19421
rect 12423 19319 12457 19353
rect 12423 19251 12457 19285
rect 12423 19183 12457 19217
rect 12423 19115 12457 19149
rect 12423 19047 12457 19081
rect 12423 18979 12457 19013
rect 12423 18911 12457 18945
rect 12423 18843 12457 18877
rect 12423 18775 12457 18809
rect 12423 18707 12457 18741
rect 12423 18639 12457 18673
rect 12423 18571 12457 18605
rect 12423 18503 12457 18537
rect 12423 18435 12457 18469
rect 12423 18367 12457 18401
rect 12423 18299 12457 18333
rect 12423 18231 12457 18265
rect 12423 18163 12457 18197
rect 12423 18095 12457 18129
rect 12423 18027 12457 18061
rect 12423 17959 12457 17993
rect 12423 17891 12457 17925
rect 12423 17823 12457 17857
rect 12423 17755 12457 17789
rect 12423 17687 12457 17721
rect 12423 17619 12457 17653
rect 12423 17551 12457 17585
rect 12423 17483 12457 17517
rect 12423 17415 12457 17449
rect 12423 17347 12457 17381
rect 12423 17279 12457 17313
rect 12423 17211 12457 17245
rect 12423 17143 12457 17177
rect 12423 17075 12457 17109
rect 12423 17007 12457 17041
rect 12423 16939 12457 16973
rect 12423 16871 12457 16905
rect 12423 16803 12457 16837
rect 12423 16735 12457 16769
rect 12423 16667 12457 16701
rect 12423 16599 12457 16633
rect 12423 16531 12457 16565
rect 12423 16463 12457 16497
rect 12423 16395 12457 16429
rect 12423 16327 12457 16361
rect 12423 16259 12457 16293
rect 12423 16191 12457 16225
rect 12423 16123 12457 16157
rect 12423 16055 12457 16089
rect 12423 15987 12457 16021
rect 12423 15919 12457 15953
rect 12423 15851 12457 15885
rect 12423 15783 12457 15817
rect 12423 15715 12457 15749
rect 12423 15647 12457 15681
rect 12423 15579 12457 15613
rect 12423 15511 12457 15545
rect 12423 15443 12457 15477
rect 12423 15375 12457 15409
rect 12423 15307 12457 15341
rect 12423 15239 12457 15273
rect 463 15163 497 15197
rect 531 15163 565 15197
rect 599 15163 633 15197
rect 667 15163 701 15197
rect 735 15163 769 15197
rect 803 15163 837 15197
rect 871 15163 905 15197
rect 939 15163 973 15197
rect 1007 15163 1041 15197
rect 1075 15163 1109 15197
rect 1143 15163 1177 15197
rect 1211 15163 1245 15197
rect 1279 15163 1313 15197
rect 1347 15163 1381 15197
rect 1415 15163 1449 15197
rect 1483 15163 1517 15197
rect 1551 15163 1585 15197
rect 1619 15163 1653 15197
rect 1687 15163 1721 15197
rect 1755 15163 1789 15197
rect 1823 15163 1857 15197
rect 1891 15163 1925 15197
rect 1959 15163 1993 15197
rect 2027 15163 2061 15197
rect 2095 15163 2129 15197
rect 2163 15163 2197 15197
rect 2231 15163 2265 15197
rect 2299 15163 2333 15197
rect 2367 15163 2401 15197
rect 2435 15163 2469 15197
rect 2503 15163 2537 15197
rect 2571 15163 2605 15197
rect 2639 15163 2673 15197
rect 2707 15163 2741 15197
rect 2775 15163 2809 15197
rect 2843 15163 2877 15197
rect 2911 15163 2945 15197
rect 2979 15163 3013 15197
rect 3047 15163 3081 15197
rect 3115 15163 3149 15197
rect 3183 15163 3217 15197
rect 3251 15163 3285 15197
rect 3319 15163 3353 15197
rect 3387 15163 3421 15197
rect 3455 15163 3489 15197
rect 3523 15163 3557 15197
rect 3591 15163 3625 15197
rect 3659 15163 3693 15197
rect 3727 15163 3761 15197
rect 3795 15163 3829 15197
rect 3863 15163 3897 15197
rect 3931 15163 3965 15197
rect 3999 15163 4033 15197
rect 4067 15163 4101 15197
rect 4135 15163 4169 15197
rect 4203 15163 4237 15197
rect 4271 15163 4305 15197
rect 4339 15163 4373 15197
rect 4407 15163 4441 15197
rect 4475 15163 4509 15197
rect 4543 15163 4577 15197
rect 4611 15163 4645 15197
rect 4679 15163 4713 15197
rect 4747 15163 4781 15197
rect 4815 15163 4849 15197
rect 4883 15163 4917 15197
rect 4951 15163 4985 15197
rect 5019 15163 5053 15197
rect 5087 15163 5121 15197
rect 5155 15163 5189 15197
rect 5223 15163 5257 15197
rect 5291 15163 5325 15197
rect 5359 15163 5393 15197
rect 5427 15163 5461 15197
rect 5495 15163 5529 15197
rect 5563 15163 5597 15197
rect 5631 15163 5665 15197
rect 5699 15163 5733 15197
rect 5767 15163 5801 15197
rect 5835 15163 5869 15197
rect 5903 15163 5937 15197
rect 5971 15163 6005 15197
rect 6039 15163 6073 15197
rect 6107 15163 6141 15197
rect 6175 15163 6209 15197
rect 6243 15163 6277 15197
rect 6311 15163 6345 15197
rect 6379 15163 6413 15197
rect 6447 15163 6481 15197
rect 6515 15163 6549 15197
rect 6583 15163 6617 15197
rect 6651 15163 6685 15197
rect 6719 15163 6753 15197
rect 6787 15163 6821 15197
rect 6855 15163 6889 15197
rect 6923 15163 6957 15197
rect 6991 15163 7025 15197
rect 7059 15163 7093 15197
rect 7127 15163 7161 15197
rect 7195 15163 7229 15197
rect 7263 15163 7297 15197
rect 7331 15163 7365 15197
rect 7399 15163 7433 15197
rect 7467 15163 7501 15197
rect 7535 15163 7569 15197
rect 7603 15163 7637 15197
rect 7671 15163 7705 15197
rect 7739 15163 7773 15197
rect 7807 15163 7841 15197
rect 7875 15163 7909 15197
rect 7943 15163 7977 15197
rect 8011 15163 8045 15197
rect 8079 15163 8113 15197
rect 8147 15163 8181 15197
rect 8215 15163 8249 15197
rect 8283 15163 8317 15197
rect 8351 15163 8385 15197
rect 8419 15163 8453 15197
rect 8487 15163 8521 15197
rect 8555 15163 8589 15197
rect 8623 15163 8657 15197
rect 8691 15163 8725 15197
rect 8759 15163 8793 15197
rect 8827 15163 8861 15197
rect 8895 15163 8929 15197
rect 8963 15163 8997 15197
rect 9031 15163 9065 15197
rect 9099 15163 9133 15197
rect 9167 15163 9201 15197
rect 9235 15163 9269 15197
rect 9303 15163 9337 15197
rect 9371 15163 9405 15197
rect 9439 15163 9473 15197
rect 9507 15163 9541 15197
rect 9575 15163 9609 15197
rect 9643 15163 9677 15197
rect 9711 15163 9745 15197
rect 9779 15163 9813 15197
rect 9847 15163 9881 15197
rect 9915 15163 9949 15197
rect 9983 15163 10017 15197
rect 10051 15163 10085 15197
rect 10119 15163 10153 15197
rect 10187 15163 10221 15197
rect 10255 15163 10289 15197
rect 10323 15163 10357 15197
rect 10391 15163 10425 15197
rect 10459 15163 10493 15197
rect 10527 15163 10561 15197
rect 10595 15163 10629 15197
rect 10663 15163 10697 15197
rect 10731 15163 10765 15197
rect 10799 15163 10833 15197
rect 10867 15163 10901 15197
rect 10935 15163 10969 15197
rect 11003 15163 11037 15197
rect 11071 15163 11105 15197
rect 11139 15163 11173 15197
rect 11207 15163 11241 15197
rect 11275 15163 11309 15197
rect 11343 15163 11377 15197
rect 11411 15163 11445 15197
rect 11479 15163 11513 15197
rect 11547 15163 11581 15197
rect 11615 15163 11649 15197
rect 11683 15163 11717 15197
rect 11751 15163 11785 15197
rect 11819 15163 11853 15197
rect 11887 15163 11921 15197
rect 11955 15163 11989 15197
rect 12023 15163 12057 15197
rect 12091 15163 12125 15197
rect 12159 15163 12193 15197
rect 12227 15163 12261 15197
rect 12295 15163 12329 15197
rect 12363 15163 12397 15197
<< locali >>
rect 403 21787 540 21817
rect 437 21783 540 21787
rect 574 21783 608 21817
rect 642 21783 676 21817
rect 710 21783 744 21817
rect 778 21783 812 21817
rect 846 21783 880 21817
rect 914 21783 948 21817
rect 982 21783 1016 21817
rect 1050 21783 1084 21817
rect 1118 21783 1152 21817
rect 1186 21783 1220 21817
rect 1254 21783 1288 21817
rect 1322 21783 1356 21817
rect 1390 21783 1424 21817
rect 1458 21783 1492 21817
rect 1526 21783 1560 21817
rect 1594 21783 1628 21817
rect 1662 21783 1696 21817
rect 1730 21783 1764 21817
rect 1798 21783 1832 21817
rect 1866 21783 1900 21817
rect 1934 21783 1968 21817
rect 2002 21783 2036 21817
rect 2070 21783 2104 21817
rect 2138 21783 2172 21817
rect 2206 21783 2240 21817
rect 2274 21783 2308 21817
rect 2342 21783 2376 21817
rect 2410 21783 2444 21817
rect 2478 21783 2512 21817
rect 2546 21783 2580 21817
rect 2614 21783 2648 21817
rect 2682 21783 2716 21817
rect 2750 21783 2784 21817
rect 2818 21783 2852 21817
rect 2886 21783 2920 21817
rect 2954 21783 2988 21817
rect 3022 21783 3056 21817
rect 3090 21783 3124 21817
rect 3158 21783 3192 21817
rect 3226 21783 3260 21817
rect 3294 21783 3328 21817
rect 3362 21783 3396 21817
rect 3430 21783 3464 21817
rect 3498 21783 3532 21817
rect 3566 21783 3600 21817
rect 3634 21783 3668 21817
rect 3702 21783 3736 21817
rect 3770 21783 3804 21817
rect 3838 21783 3872 21817
rect 3906 21783 3940 21817
rect 3974 21783 4008 21817
rect 4042 21783 4076 21817
rect 4110 21783 4144 21817
rect 4178 21783 4212 21817
rect 4246 21783 4280 21817
rect 4314 21783 4348 21817
rect 4382 21783 4416 21817
rect 4450 21783 4484 21817
rect 4518 21783 4552 21817
rect 4586 21783 4620 21817
rect 4654 21783 4688 21817
rect 4722 21783 4756 21817
rect 4790 21783 4824 21817
rect 4858 21783 4892 21817
rect 4926 21783 4960 21817
rect 4994 21783 5028 21817
rect 5062 21783 5096 21817
rect 5130 21783 5164 21817
rect 5198 21783 5232 21817
rect 5266 21783 5300 21817
rect 5334 21783 5368 21817
rect 5402 21783 5436 21817
rect 5470 21783 5504 21817
rect 5538 21783 5572 21817
rect 5606 21783 5640 21817
rect 5674 21783 5708 21817
rect 5742 21783 5776 21817
rect 5810 21783 5844 21817
rect 5878 21783 5912 21817
rect 5946 21783 5980 21817
rect 6014 21783 6048 21817
rect 6082 21783 6116 21817
rect 6150 21783 6184 21817
rect 6218 21783 6252 21817
rect 6286 21783 6320 21817
rect 6354 21783 6388 21817
rect 6422 21783 6456 21817
rect 6490 21783 6524 21817
rect 6558 21783 6592 21817
rect 6626 21783 6660 21817
rect 6694 21783 6728 21817
rect 6762 21783 6796 21817
rect 6830 21783 6864 21817
rect 6898 21783 6932 21817
rect 6966 21783 7000 21817
rect 7034 21783 7068 21817
rect 7102 21783 7136 21817
rect 7170 21783 7204 21817
rect 7238 21783 7272 21817
rect 7306 21783 7340 21817
rect 7374 21783 7408 21817
rect 7442 21783 7476 21817
rect 7510 21783 7544 21817
rect 7578 21783 7612 21817
rect 7646 21783 7680 21817
rect 7714 21783 7748 21817
rect 7782 21783 7816 21817
rect 7850 21783 7884 21817
rect 7918 21783 7952 21817
rect 7986 21783 8020 21817
rect 8054 21783 8088 21817
rect 8122 21783 8156 21817
rect 8190 21783 8224 21817
rect 8258 21783 8292 21817
rect 8326 21783 8360 21817
rect 8394 21783 8428 21817
rect 8462 21783 8496 21817
rect 8530 21783 8564 21817
rect 8598 21783 8632 21817
rect 8666 21783 8700 21817
rect 8734 21783 8768 21817
rect 8802 21783 8836 21817
rect 8870 21783 8904 21817
rect 8938 21783 8972 21817
rect 9006 21783 9040 21817
rect 9074 21783 9108 21817
rect 9142 21783 9176 21817
rect 9210 21783 9244 21817
rect 9278 21783 9312 21817
rect 9346 21783 9380 21817
rect 9414 21783 9448 21817
rect 9482 21783 9516 21817
rect 9550 21783 9584 21817
rect 9618 21783 9652 21817
rect 9686 21783 9720 21817
rect 9754 21783 9788 21817
rect 9822 21783 9856 21817
rect 9890 21783 9924 21817
rect 9958 21783 9992 21817
rect 10026 21783 10060 21817
rect 10094 21783 10128 21817
rect 10162 21783 10196 21817
rect 10230 21783 10264 21817
rect 10298 21783 10332 21817
rect 10366 21783 10400 21817
rect 10434 21783 10468 21817
rect 10502 21783 10536 21817
rect 10570 21783 10604 21817
rect 10638 21783 10672 21817
rect 10706 21783 10740 21817
rect 10774 21783 10808 21817
rect 10842 21783 10876 21817
rect 10910 21783 10944 21817
rect 10978 21783 11012 21817
rect 11046 21783 11080 21817
rect 11114 21783 11148 21817
rect 11182 21783 11216 21817
rect 11250 21783 11284 21817
rect 11318 21783 11352 21817
rect 11386 21783 11420 21817
rect 11454 21783 11488 21817
rect 11522 21783 11556 21817
rect 11590 21783 11624 21817
rect 11658 21783 11692 21817
rect 11726 21783 11760 21817
rect 11794 21783 11828 21817
rect 11862 21783 11896 21817
rect 11930 21783 11964 21817
rect 11998 21783 12032 21817
rect 12066 21783 12100 21817
rect 12134 21783 12168 21817
rect 12202 21783 12236 21817
rect 12270 21783 12304 21817
rect 12338 21783 12457 21817
rect 12480 21783 12510 21817
rect 403 21719 437 21753
rect 403 21651 437 21685
rect 403 21583 437 21617
rect 403 21515 437 21549
rect 403 21447 437 21481
rect 12423 21733 12457 21783
rect 12423 21665 12457 21699
rect 12423 21597 12457 21631
rect 12423 21529 12457 21563
rect 403 21379 437 21413
rect 1030 21442 1280 21470
rect 1064 21408 1075 21442
rect 1136 21408 1143 21442
rect 1208 21408 1211 21442
rect 1245 21408 1246 21442
rect 1030 21380 1280 21408
rect 7010 21437 7280 21470
rect 7010 21403 7020 21437
rect 7054 21403 7055 21437
rect 7089 21403 7092 21437
rect 7157 21403 7164 21437
rect 7225 21403 7236 21437
rect 7270 21403 7280 21437
rect 7010 21370 7280 21403
rect 12423 21461 12457 21495
rect 12423 21393 12457 21427
rect 403 21311 437 21345
rect 403 21243 437 21277
rect 403 21175 437 21209
rect 403 21107 437 21141
rect 403 21039 437 21073
rect 403 20971 437 21005
rect 403 20903 437 20937
rect 403 20835 437 20869
rect 403 20767 437 20801
rect 403 20699 437 20733
rect 403 20631 437 20665
rect 403 20563 437 20597
rect 403 20495 437 20529
rect 403 20427 437 20461
rect 403 20359 437 20393
rect 403 20291 437 20325
rect 403 20223 437 20257
rect 403 20155 437 20189
rect 403 20087 437 20121
rect 403 20019 437 20053
rect 403 19951 437 19985
rect 403 19883 437 19917
rect 403 19815 437 19849
rect 403 19747 437 19781
rect 403 19679 437 19713
rect 403 19611 437 19645
rect 403 19543 437 19577
rect 403 19475 437 19509
rect 403 19407 437 19441
rect 403 19339 437 19373
rect 403 19271 437 19305
rect 403 19203 437 19237
rect 403 19135 437 19169
rect 403 19067 437 19101
rect 403 18999 437 19033
rect 403 18931 437 18965
rect 403 18863 437 18897
rect 403 18795 437 18829
rect 403 18727 437 18761
rect 403 18659 437 18693
rect 403 18591 437 18625
rect 403 18523 437 18557
rect 403 18455 437 18489
rect 403 18387 437 18421
rect 403 18319 437 18353
rect 403 18251 437 18285
rect 403 18183 437 18217
rect 403 18115 437 18149
rect 403 18047 437 18081
rect 403 17979 437 18013
rect 403 17911 437 17945
rect 403 17843 437 17877
rect 403 17775 437 17809
rect 403 17707 437 17741
rect 403 17639 437 17673
rect 403 17571 437 17605
rect 403 17503 437 17537
rect 403 17435 437 17469
rect 403 17367 437 17401
rect 403 17299 437 17333
rect 403 17231 437 17265
rect 403 17163 437 17197
rect 403 17095 437 17129
rect 403 17027 437 17061
rect 403 16959 437 16993
rect 403 16891 437 16925
rect 403 16823 437 16857
rect 403 16755 437 16789
rect 403 16687 437 16721
rect 403 16619 437 16653
rect 403 16551 437 16585
rect 403 16483 437 16517
rect 403 16415 437 16449
rect 403 16347 437 16381
rect 403 16279 437 16313
rect 403 16211 437 16245
rect 403 16143 437 16177
rect 403 16075 437 16109
rect 403 16007 437 16041
rect 403 15939 437 15973
rect 403 15871 437 15905
rect 403 15803 437 15837
rect 403 15735 437 15769
rect 403 15667 437 15701
rect 403 15599 437 15633
rect 403 15531 437 15565
rect 403 15463 437 15497
rect 403 15395 437 15429
rect 403 15327 437 15361
rect 403 15259 437 15293
rect 403 15197 437 15225
rect 12423 21325 12457 21359
rect 12423 21257 12457 21291
rect 12423 21189 12457 21223
rect 12423 21121 12457 21155
rect 12423 21053 12457 21087
rect 12423 20985 12457 21019
rect 12423 20917 12457 20951
rect 12423 20849 12457 20883
rect 12423 20781 12457 20815
rect 12423 20713 12457 20747
rect 12423 20645 12457 20679
rect 12423 20577 12457 20611
rect 12423 20509 12457 20543
rect 12423 20441 12457 20475
rect 12423 20373 12457 20407
rect 12423 20305 12457 20339
rect 12423 20237 12457 20271
rect 12423 20169 12457 20203
rect 12423 20101 12457 20135
rect 12423 20033 12457 20067
rect 12423 19965 12457 19999
rect 12423 19897 12457 19931
rect 12423 19829 12457 19863
rect 12423 19761 12457 19795
rect 12423 19693 12457 19727
rect 12423 19625 12457 19659
rect 12423 19557 12457 19591
rect 12423 19489 12457 19523
rect 12423 19421 12457 19455
rect 12423 19353 12457 19387
rect 12423 19285 12457 19319
rect 12423 19217 12457 19251
rect 12423 19149 12457 19183
rect 12423 19081 12457 19115
rect 12423 19013 12457 19047
rect 12423 18945 12457 18979
rect 12423 18877 12457 18911
rect 12423 18809 12457 18843
rect 12423 18741 12457 18775
rect 12423 18673 12457 18707
rect 12423 18605 12457 18639
rect 12423 18537 12457 18571
rect 12423 18469 12457 18503
rect 12423 18401 12457 18435
rect 12423 18333 12457 18367
rect 12423 18265 12457 18299
rect 12423 18197 12457 18231
rect 12423 18129 12457 18163
rect 12423 18061 12457 18095
rect 12423 17993 12457 18027
rect 12423 17925 12457 17959
rect 12423 17857 12457 17891
rect 12423 17789 12457 17823
rect 12423 17721 12457 17755
rect 12423 17653 12457 17687
rect 12423 17585 12457 17619
rect 12423 17517 12457 17551
rect 12423 17449 12457 17483
rect 12423 17381 12457 17415
rect 12423 17313 12457 17347
rect 12423 17245 12457 17279
rect 12423 17177 12457 17211
rect 12423 17109 12457 17143
rect 12423 17041 12457 17075
rect 12423 16973 12457 17007
rect 12423 16905 12457 16939
rect 12423 16837 12457 16871
rect 12423 16769 12457 16803
rect 12423 16701 12457 16735
rect 12423 16633 12457 16667
rect 12423 16565 12457 16599
rect 12423 16497 12457 16531
rect 12423 16429 12457 16463
rect 12423 16361 12457 16395
rect 12423 16293 12457 16327
rect 12423 16225 12457 16259
rect 12423 16157 12457 16191
rect 12423 16089 12457 16123
rect 12423 16021 12457 16055
rect 12423 15953 12457 15987
rect 12423 15885 12457 15919
rect 12423 15817 12457 15851
rect 12423 15749 12457 15783
rect 12423 15681 12457 15715
rect 12423 15613 12457 15647
rect 12423 15545 12457 15579
rect 12423 15477 12457 15511
rect 12423 15409 12457 15443
rect 12423 15341 12457 15375
rect 12423 15273 12457 15307
rect 12423 15197 12457 15239
rect 403 15163 463 15197
rect 497 15163 531 15197
rect 565 15163 599 15197
rect 633 15163 667 15197
rect 701 15163 735 15197
rect 769 15163 803 15197
rect 837 15163 871 15197
rect 905 15163 939 15197
rect 973 15163 1007 15197
rect 1041 15163 1075 15197
rect 1109 15163 1143 15197
rect 1177 15163 1211 15197
rect 1245 15163 1279 15197
rect 1313 15163 1347 15197
rect 1381 15163 1415 15197
rect 1449 15163 1483 15197
rect 1517 15163 1551 15197
rect 1585 15163 1619 15197
rect 1653 15163 1687 15197
rect 1721 15163 1755 15197
rect 1789 15163 1823 15197
rect 1857 15163 1891 15197
rect 1925 15163 1959 15197
rect 1993 15163 2027 15197
rect 2061 15163 2095 15197
rect 2129 15163 2163 15197
rect 2197 15163 2231 15197
rect 2265 15163 2299 15197
rect 2333 15163 2367 15197
rect 2401 15163 2435 15197
rect 2469 15163 2503 15197
rect 2537 15163 2571 15197
rect 2605 15163 2639 15197
rect 2673 15163 2707 15197
rect 2741 15163 2775 15197
rect 2809 15163 2843 15197
rect 2877 15163 2911 15197
rect 2945 15163 2979 15197
rect 3013 15163 3047 15197
rect 3081 15163 3115 15197
rect 3149 15163 3183 15197
rect 3217 15163 3251 15197
rect 3285 15163 3319 15197
rect 3353 15163 3387 15197
rect 3421 15163 3455 15197
rect 3489 15163 3523 15197
rect 3557 15163 3591 15197
rect 3625 15163 3659 15197
rect 3693 15163 3727 15197
rect 3761 15163 3795 15197
rect 3829 15163 3863 15197
rect 3897 15163 3931 15197
rect 3965 15163 3999 15197
rect 4033 15163 4067 15197
rect 4101 15163 4135 15197
rect 4169 15163 4203 15197
rect 4237 15163 4271 15197
rect 4305 15163 4339 15197
rect 4373 15163 4407 15197
rect 4441 15163 4475 15197
rect 4509 15163 4543 15197
rect 4577 15163 4611 15197
rect 4645 15163 4679 15197
rect 4713 15163 4747 15197
rect 4781 15163 4815 15197
rect 4849 15163 4883 15197
rect 4917 15163 4951 15197
rect 4985 15163 5019 15197
rect 5053 15163 5087 15197
rect 5121 15163 5155 15197
rect 5189 15163 5223 15197
rect 5257 15163 5291 15197
rect 5325 15163 5359 15197
rect 5393 15163 5427 15197
rect 5461 15163 5495 15197
rect 5529 15163 5563 15197
rect 5597 15163 5631 15197
rect 5665 15163 5699 15197
rect 5733 15163 5767 15197
rect 5801 15163 5835 15197
rect 5869 15163 5903 15197
rect 5937 15163 5971 15197
rect 6005 15163 6039 15197
rect 6073 15163 6107 15197
rect 6141 15163 6175 15197
rect 6209 15163 6243 15197
rect 6277 15163 6311 15197
rect 6345 15163 6379 15197
rect 6413 15163 6447 15197
rect 6481 15163 6515 15197
rect 6549 15163 6583 15197
rect 6617 15163 6651 15197
rect 6685 15163 6719 15197
rect 6753 15163 6787 15197
rect 6821 15163 6855 15197
rect 6889 15163 6923 15197
rect 6957 15163 6991 15197
rect 7025 15163 7059 15197
rect 7093 15163 7127 15197
rect 7161 15163 7195 15197
rect 7229 15163 7263 15197
rect 7297 15163 7331 15197
rect 7365 15163 7399 15197
rect 7433 15163 7467 15197
rect 7501 15163 7535 15197
rect 7569 15163 7603 15197
rect 7637 15163 7671 15197
rect 7705 15163 7739 15197
rect 7773 15163 7807 15197
rect 7841 15163 7875 15197
rect 7909 15163 7943 15197
rect 7977 15163 8011 15197
rect 8045 15163 8079 15197
rect 8113 15163 8147 15197
rect 8181 15163 8215 15197
rect 8249 15163 8283 15197
rect 8317 15163 8351 15197
rect 8385 15163 8419 15197
rect 8453 15163 8487 15197
rect 8521 15163 8555 15197
rect 8589 15163 8623 15197
rect 8657 15163 8691 15197
rect 8725 15163 8759 15197
rect 8793 15163 8827 15197
rect 8861 15163 8895 15197
rect 8929 15163 8963 15197
rect 8997 15163 9031 15197
rect 9065 15163 9099 15197
rect 9133 15163 9167 15197
rect 9201 15163 9235 15197
rect 9269 15163 9303 15197
rect 9337 15163 9371 15197
rect 9405 15163 9439 15197
rect 9473 15163 9507 15197
rect 9541 15163 9575 15197
rect 9609 15163 9643 15197
rect 9677 15163 9711 15197
rect 9745 15163 9779 15197
rect 9813 15163 9847 15197
rect 9881 15163 9915 15197
rect 9949 15163 9983 15197
rect 10017 15163 10051 15197
rect 10085 15163 10119 15197
rect 10153 15163 10187 15197
rect 10221 15163 10255 15197
rect 10289 15163 10323 15197
rect 10357 15163 10391 15197
rect 10425 15163 10459 15197
rect 10493 15163 10527 15197
rect 10561 15163 10595 15197
rect 10629 15163 10663 15197
rect 10697 15163 10731 15197
rect 10765 15163 10799 15197
rect 10833 15163 10867 15197
rect 10901 15163 10935 15197
rect 10969 15163 11003 15197
rect 11037 15163 11071 15197
rect 11105 15163 11139 15197
rect 11173 15163 11207 15197
rect 11241 15163 11275 15197
rect 11309 15163 11343 15197
rect 11377 15163 11411 15197
rect 11445 15163 11479 15197
rect 11513 15163 11547 15197
rect 11581 15163 11615 15197
rect 11649 15163 11683 15197
rect 11717 15163 11751 15197
rect 11785 15163 11819 15197
rect 11853 15163 11887 15197
rect 11921 15163 11955 15197
rect 11989 15163 12023 15197
rect 12057 15163 12091 15197
rect 12125 15163 12159 15197
rect 12193 15163 12227 15197
rect 12261 15163 12295 15197
rect 12329 15163 12363 15197
rect 12397 15163 12457 15197
rect 383 13183 458 13217
rect 492 13183 526 13217
rect 560 13183 594 13217
rect 628 13183 662 13217
rect 696 13183 730 13217
rect 764 13183 798 13217
rect 832 13183 866 13217
rect 900 13183 934 13217
rect 968 13183 1002 13217
rect 1036 13183 1070 13217
rect 1104 13183 1138 13217
rect 1172 13183 1206 13217
rect 1240 13183 1274 13217
rect 1308 13183 1342 13217
rect 1376 13183 1410 13217
rect 1444 13183 1478 13217
rect 1512 13183 1546 13217
rect 1580 13183 1614 13217
rect 1648 13183 1682 13217
rect 1716 13183 1750 13217
rect 1784 13183 1818 13217
rect 1852 13183 1886 13217
rect 1920 13183 1954 13217
rect 1988 13183 2022 13217
rect 2056 13183 2090 13217
rect 2124 13183 2158 13217
rect 2192 13183 2226 13217
rect 2260 13183 2294 13217
rect 2328 13183 2362 13217
rect 2396 13183 2430 13217
rect 2464 13183 2498 13217
rect 2532 13183 2566 13217
rect 2600 13183 2634 13217
rect 2668 13183 2702 13217
rect 2736 13183 2770 13217
rect 2804 13183 2838 13217
rect 2872 13183 2906 13217
rect 2940 13183 2974 13217
rect 3008 13183 3042 13217
rect 3076 13183 3110 13217
rect 3144 13183 3178 13217
rect 3212 13183 3246 13217
rect 3280 13183 3314 13217
rect 3348 13183 3382 13217
rect 3416 13183 3450 13217
rect 3484 13183 3518 13217
rect 3552 13183 3586 13217
rect 3620 13183 3654 13217
rect 3688 13183 3722 13217
rect 3756 13183 3790 13217
rect 3824 13183 3858 13217
rect 3892 13183 3926 13217
rect 3960 13183 3994 13217
rect 4028 13183 4062 13217
rect 4096 13183 4130 13217
rect 4164 13183 4198 13217
rect 4232 13183 4266 13217
rect 4300 13183 4334 13217
rect 4368 13183 4402 13217
rect 4436 13183 4470 13217
rect 4504 13183 4538 13217
rect 4572 13183 4606 13217
rect 4640 13183 4674 13217
rect 4708 13183 4742 13217
rect 4776 13183 4810 13217
rect 4844 13183 4878 13217
rect 4912 13183 4946 13217
rect 4980 13183 5014 13217
rect 5048 13183 5082 13217
rect 5116 13183 5150 13217
rect 5184 13183 5218 13217
rect 5252 13183 5286 13217
rect 5320 13183 5354 13217
rect 5388 13183 5422 13217
rect 5456 13183 5490 13217
rect 5524 13183 5558 13217
rect 5592 13183 5626 13217
rect 5660 13183 5694 13217
rect 5728 13183 5762 13217
rect 5796 13183 5830 13217
rect 5864 13183 5898 13217
rect 5932 13183 5966 13217
rect 6000 13183 6034 13217
rect 6068 13183 6102 13217
rect 6136 13183 6170 13217
rect 6204 13183 6238 13217
rect 6272 13183 6306 13217
rect 6340 13183 6374 13217
rect 6408 13183 6442 13217
rect 6476 13183 6510 13217
rect 6544 13183 6578 13217
rect 6612 13183 6646 13217
rect 6680 13183 6714 13217
rect 6748 13183 6782 13217
rect 6816 13183 6850 13217
rect 6884 13183 6918 13217
rect 6952 13183 6986 13217
rect 7020 13183 7054 13217
rect 7088 13183 7122 13217
rect 7156 13183 7190 13217
rect 7224 13183 7258 13217
rect 7292 13183 7326 13217
rect 7360 13183 7394 13217
rect 7428 13183 7462 13217
rect 7496 13183 7530 13217
rect 7564 13183 7598 13217
rect 7632 13183 7666 13217
rect 7700 13183 7734 13217
rect 7768 13183 7802 13217
rect 7836 13183 7870 13217
rect 7904 13183 7938 13217
rect 7972 13183 8006 13217
rect 8040 13183 8074 13217
rect 8108 13183 8142 13217
rect 8176 13183 8210 13217
rect 8244 13183 8278 13217
rect 8312 13183 8346 13217
rect 8380 13183 8414 13217
rect 8448 13183 8482 13217
rect 8516 13183 8550 13217
rect 8584 13183 8618 13217
rect 8652 13183 8686 13217
rect 8720 13183 8754 13217
rect 8788 13183 8822 13217
rect 8856 13183 8890 13217
rect 8924 13183 8958 13217
rect 8992 13183 9026 13217
rect 9060 13183 9094 13217
rect 9128 13183 9162 13217
rect 9196 13183 9230 13217
rect 9264 13183 9384 13217
rect 9418 13183 9452 13217
rect 9486 13183 9520 13217
rect 9554 13183 9588 13217
rect 9622 13183 9656 13217
rect 9690 13183 9724 13217
rect 9758 13183 9792 13217
rect 9826 13183 9860 13217
rect 9894 13183 9928 13217
rect 9962 13183 9996 13217
rect 10030 13183 10064 13217
rect 10098 13183 10132 13217
rect 10166 13183 10200 13217
rect 10234 13183 10268 13217
rect 10302 13183 10336 13217
rect 10370 13183 10404 13217
rect 10438 13183 10472 13217
rect 10506 13183 10540 13217
rect 10574 13183 10608 13217
rect 10642 13183 10676 13217
rect 10710 13183 10744 13217
rect 10778 13183 10812 13217
rect 10846 13183 10880 13217
rect 10914 13183 10948 13217
rect 10982 13183 11016 13217
rect 11050 13183 11084 13217
rect 11118 13183 11152 13217
rect 11186 13183 11220 13217
rect 11254 13183 11288 13217
rect 11322 13183 11356 13217
rect 11390 13183 11424 13217
rect 11458 13183 11492 13217
rect 11526 13183 11607 13217
rect 383 13135 417 13183
rect 383 13067 417 13101
rect 383 12999 417 13033
rect 383 12931 417 12965
rect 383 12863 417 12897
rect 383 12795 417 12829
rect 383 12727 417 12761
rect 383 12659 417 12693
rect 383 12591 417 12625
rect 383 12523 417 12557
rect 383 12455 417 12489
rect 383 12387 417 12421
rect 11573 13137 11607 13183
rect 11573 13069 11607 13103
rect 11573 13001 11607 13035
rect 11573 12933 11607 12967
rect 11573 12865 11607 12899
rect 11573 12797 11607 12831
rect 11573 12729 11607 12763
rect 11573 12661 11607 12695
rect 11573 12593 11607 12627
rect 11573 12525 11607 12559
rect 11573 12457 11607 12491
rect 383 12319 417 12353
rect 383 12251 417 12285
rect 2690 12347 2790 12396
rect 2690 12313 2723 12347
rect 2757 12313 2790 12347
rect 2690 12264 2790 12313
rect 2870 12347 2970 12396
rect 11573 12389 11607 12423
rect 2870 12313 2903 12347
rect 2937 12313 2970 12347
rect 2870 12264 2970 12313
rect 5590 12337 5690 12386
rect 5590 12303 5623 12337
rect 5657 12303 5690 12337
rect 5590 12254 5690 12303
rect 5770 12337 5870 12386
rect 5770 12303 5803 12337
rect 5837 12303 5870 12337
rect 5770 12254 5870 12303
rect 11573 12321 11607 12355
rect 383 12183 417 12217
rect 383 12115 417 12149
rect 383 12047 417 12081
rect 383 11979 417 12013
rect 383 11911 417 11945
rect 383 11843 417 11877
rect 383 11775 417 11809
rect 383 11707 417 11741
rect 383 11639 417 11673
rect 383 11571 417 11605
rect 383 11503 417 11537
rect 383 11435 417 11469
rect 383 11367 417 11401
rect 383 11299 417 11333
rect 383 11231 417 11265
rect 383 11163 417 11197
rect 383 11095 417 11129
rect 383 11027 417 11061
rect 383 10959 417 10993
rect 11573 12253 11607 12287
rect 11573 12185 11607 12219
rect 11573 12117 11607 12151
rect 11573 12049 11607 12083
rect 11573 11981 11607 12015
rect 11573 11913 11607 11947
rect 11573 11845 11607 11879
rect 11573 11777 11607 11811
rect 11573 11709 11607 11743
rect 11573 11641 11607 11675
rect 11573 11573 11607 11607
rect 11573 11505 11607 11539
rect 11573 11437 11607 11471
rect 11573 11369 11607 11403
rect 11573 11301 11607 11335
rect 11573 11233 11607 11267
rect 11573 11165 11607 11199
rect 11573 11097 11607 11131
rect 11573 11017 11607 11063
rect 11573 10983 11644 11017
rect 11678 10983 11712 11017
rect 11746 10983 11780 11017
rect 11814 10983 11848 11017
rect 11882 10983 11916 11017
rect 11950 10983 11984 11017
rect 12018 10983 12052 11017
rect 12086 10983 12120 11017
rect 12154 10983 12188 11017
rect 12222 10983 12256 11017
rect 12290 10983 12324 11017
rect 12358 10983 12392 11017
rect 12426 10983 12460 11017
rect 12494 10983 12528 11017
rect 12562 10983 12596 11017
rect 12630 10983 12664 11017
rect 12698 10983 12732 11017
rect 12766 10983 12800 11017
rect 12834 10983 12868 11017
rect 12902 10983 12936 11017
rect 12970 10983 13004 11017
rect 13038 10983 13072 11017
rect 13106 10983 13140 11017
rect 13174 10983 13208 11017
rect 13242 10983 13276 11017
rect 13310 10983 13344 11017
rect 13378 10983 13412 11017
rect 13446 10983 13480 11017
rect 13514 10983 13548 11017
rect 13582 10983 13616 11017
rect 13650 10983 13684 11017
rect 13718 10983 13752 11017
rect 13786 10983 13820 11017
rect 13854 10983 13888 11017
rect 13922 10983 13956 11017
rect 13990 10983 14024 11017
rect 14058 10983 14092 11017
rect 14126 10983 14160 11017
rect 14194 10983 14228 11017
rect 14262 10983 14296 11017
rect 14330 10983 14364 11017
rect 14398 10983 14432 11017
rect 14466 10983 14500 11017
rect 14534 10983 14568 11017
rect 14602 10983 14636 11017
rect 14670 10983 14704 11017
rect 14738 10983 14772 11017
rect 14806 10983 14840 11017
rect 14874 10983 14908 11017
rect 14942 10983 14976 11017
rect 15010 10983 15044 11017
rect 15078 10983 15112 11017
rect 15146 10983 15180 11017
rect 15214 10983 15248 11017
rect 15282 10983 15316 11017
rect 15350 10983 15384 11017
rect 15418 10983 15452 11017
rect 15486 10983 15520 11017
rect 15554 10983 15588 11017
rect 15622 10983 15656 11017
rect 15690 10983 15724 11017
rect 15758 10983 15792 11017
rect 15826 10983 15860 11017
rect 15894 10983 15928 11017
rect 15962 10983 15996 11017
rect 16030 10983 16064 11017
rect 16098 10983 16132 11017
rect 16166 10983 16200 11017
rect 16234 10983 16268 11017
rect 16302 10983 16336 11017
rect 16370 10983 16404 11017
rect 16438 10983 16472 11017
rect 16506 10983 16540 11017
rect 16574 10983 16608 11017
rect 16642 10983 16676 11017
rect 16710 10983 16744 11017
rect 16778 10983 16812 11017
rect 16846 10983 16880 11017
rect 16914 10983 16948 11017
rect 16982 10983 17016 11017
rect 17050 10983 17084 11017
rect 17118 10983 17152 11017
rect 17186 10983 17220 11017
rect 17254 10983 17288 11017
rect 17322 10983 17356 11017
rect 17390 10983 17424 11017
rect 17458 10983 17492 11017
rect 17526 10983 17560 11017
rect 17594 10983 17628 11017
rect 17662 10983 17696 11017
rect 17730 10983 17764 11017
rect 17798 10983 17832 11017
rect 17866 10983 17900 11017
rect 17934 10983 17968 11017
rect 18002 10983 18036 11017
rect 18070 10983 18104 11017
rect 18138 10983 18172 11017
rect 18206 10983 18240 11017
rect 18274 10983 18308 11017
rect 18342 10983 18376 11017
rect 18410 10983 18444 11017
rect 18478 10983 18512 11017
rect 18546 10983 18580 11017
rect 18614 10983 18648 11017
rect 18682 10983 18716 11017
rect 18750 10983 18784 11017
rect 18818 10983 18852 11017
rect 18886 10983 18920 11017
rect 18954 10983 18988 11017
rect 19022 10983 19056 11017
rect 19090 10983 19124 11017
rect 19158 10983 19192 11017
rect 19226 10983 19260 11017
rect 19294 10983 19328 11017
rect 19362 10983 19396 11017
rect 19430 10983 19464 11017
rect 19498 10983 19532 11017
rect 19566 10983 19600 11017
rect 19634 10983 19668 11017
rect 19702 10983 19736 11017
rect 19770 10983 19804 11017
rect 19838 10983 19872 11017
rect 19906 10983 19940 11017
rect 19974 10983 20008 11017
rect 20042 10983 20076 11017
rect 20110 10983 20144 11017
rect 20178 10983 20212 11017
rect 20246 10983 20280 11017
rect 20314 10983 20348 11017
rect 20382 10983 20416 11017
rect 20450 10983 20484 11017
rect 20518 10983 20552 11017
rect 20586 10983 20620 11017
rect 20654 10983 20688 11017
rect 20722 10983 20756 11017
rect 20790 10983 20824 11017
rect 20858 10983 20892 11017
rect 20926 10983 20960 11017
rect 20994 10983 21028 11017
rect 21062 10983 21096 11017
rect 21130 10983 21164 11017
rect 21198 10983 21232 11017
rect 21266 10983 21300 11017
rect 21334 10983 21368 11017
rect 21402 10983 21436 11017
rect 21470 10983 21504 11017
rect 21538 10983 21572 11017
rect 21606 10983 21640 11017
rect 21674 10983 21708 11017
rect 21742 10983 21776 11017
rect 21810 10983 21844 11017
rect 21878 10983 21912 11017
rect 21946 10983 21980 11017
rect 22014 10983 22048 11017
rect 22082 10983 22116 11017
rect 22150 10983 22184 11017
rect 22218 10983 22252 11017
rect 22286 10983 22320 11017
rect 22354 10983 22388 11017
rect 22422 10983 22497 11017
rect 383 10891 417 10925
rect 383 10823 417 10857
rect 383 10755 417 10789
rect 383 10687 417 10721
rect 383 10619 417 10653
rect 383 10551 417 10585
rect 383 10483 417 10517
rect 383 10415 417 10449
rect 22463 10947 22497 10983
rect 22463 10879 22497 10913
rect 22463 10811 22497 10845
rect 22463 10743 22497 10777
rect 22463 10675 22497 10709
rect 22463 10607 22497 10641
rect 22463 10539 22497 10573
rect 22463 10471 22497 10505
rect 383 10347 417 10381
rect 14260 10407 14420 10440
rect 14260 10373 14323 10407
rect 14357 10373 14420 10407
rect 14260 10340 14420 10373
rect 22463 10403 22497 10437
rect 383 10279 417 10313
rect 383 10211 417 10245
rect 383 10143 417 10177
rect 383 10075 417 10109
rect 383 10007 417 10041
rect 383 9939 417 9973
rect 383 9871 417 9905
rect 383 9803 417 9837
rect 383 9735 417 9769
rect 383 9667 417 9701
rect 383 9599 417 9633
rect 383 9531 417 9565
rect 383 9463 417 9497
rect 383 9395 417 9429
rect 383 9327 417 9361
rect 383 9259 417 9293
rect 383 9191 417 9225
rect 383 9123 417 9157
rect 383 9055 417 9089
rect 383 8987 417 9021
rect 383 8919 417 8953
rect 383 8851 417 8885
rect 383 8783 417 8817
rect 383 8715 417 8749
rect 383 8647 417 8681
rect 383 8579 417 8613
rect 383 8511 417 8545
rect 383 8443 417 8477
rect 383 8375 417 8409
rect 383 8307 417 8341
rect 383 8239 417 8273
rect 383 8171 417 8205
rect 383 8103 417 8137
rect 383 8035 417 8069
rect 383 7967 417 8001
rect 383 7899 417 7933
rect 383 7831 417 7865
rect 383 7763 417 7797
rect 383 7695 417 7729
rect 383 7627 417 7661
rect 383 7559 417 7593
rect 383 7491 417 7525
rect 383 7423 417 7457
rect 383 7355 417 7389
rect 383 7287 417 7321
rect 383 7219 417 7253
rect 383 7151 417 7185
rect 383 7083 417 7117
rect 383 7015 417 7049
rect 383 6947 417 6981
rect 383 6879 417 6913
rect 383 6811 417 6845
rect 383 6743 417 6777
rect 383 6675 417 6709
rect 383 6607 417 6641
rect 383 6539 417 6573
rect 383 6471 417 6505
rect 383 6403 417 6437
rect 383 6335 417 6369
rect 383 6267 417 6301
rect 383 6199 417 6233
rect 383 6131 417 6165
rect 383 6063 417 6097
rect 383 5995 417 6029
rect 383 5927 417 5961
rect 22463 10335 22497 10369
rect 22463 10267 22497 10301
rect 22463 10199 22497 10233
rect 22463 10131 22497 10165
rect 22463 10063 22497 10097
rect 22463 9995 22497 10029
rect 22463 9927 22497 9961
rect 22463 9859 22497 9893
rect 22463 9791 22497 9825
rect 22463 9723 22497 9757
rect 22463 9655 22497 9689
rect 22463 9587 22497 9621
rect 22463 9519 22497 9553
rect 22463 9451 22497 9485
rect 22463 9383 22497 9417
rect 22463 9315 22497 9349
rect 22463 9247 22497 9281
rect 22463 9179 22497 9213
rect 22463 9111 22497 9145
rect 22463 9043 22497 9077
rect 22463 8975 22497 9009
rect 22463 8907 22497 8941
rect 22463 8839 22497 8873
rect 22463 8771 22497 8805
rect 22463 8703 22497 8737
rect 22463 8635 22497 8669
rect 22463 8567 22497 8601
rect 22463 8499 22497 8533
rect 22463 8431 22497 8465
rect 22463 8363 22497 8397
rect 22463 8295 22497 8329
rect 22463 8227 22497 8261
rect 22463 8159 22497 8193
rect 22463 8091 22497 8125
rect 22463 8023 22497 8057
rect 22463 7955 22497 7989
rect 22463 7887 22497 7921
rect 22463 7819 22497 7853
rect 22463 7751 22497 7785
rect 22463 7683 22497 7717
rect 22463 7615 22497 7649
rect 22463 7547 22497 7581
rect 22463 7479 22497 7513
rect 22463 7411 22497 7445
rect 22463 7343 22497 7377
rect 22463 7275 22497 7309
rect 22463 7207 22497 7241
rect 22463 7139 22497 7173
rect 22463 7071 22497 7105
rect 22463 7003 22497 7037
rect 22463 6935 22497 6969
rect 22463 6867 22497 6901
rect 22463 6799 22497 6833
rect 22463 6731 22497 6765
rect 22463 6663 22497 6697
rect 22463 6595 22497 6629
rect 22463 6527 22497 6561
rect 22463 6459 22497 6493
rect 22463 6391 22497 6425
rect 22463 6323 22497 6357
rect 22463 6255 22497 6289
rect 22463 6187 22497 6221
rect 22463 6119 22497 6153
rect 22463 6051 22497 6085
rect 22463 5983 22497 6017
rect 383 5859 417 5893
rect 383 5791 417 5825
rect 1590 5877 1690 5926
rect 1590 5843 1623 5877
rect 1657 5843 1690 5877
rect 1590 5794 1690 5843
rect 22463 5915 22497 5949
rect 22463 5847 22497 5881
rect 383 5723 417 5757
rect 383 5655 417 5689
rect 383 5587 417 5621
rect 383 5519 417 5553
rect 383 5451 417 5485
rect 383 5383 417 5417
rect 383 5315 417 5349
rect 383 5247 417 5281
rect 383 5179 417 5213
rect 383 5111 417 5145
rect 383 5043 417 5077
rect 383 4975 417 5009
rect 383 4907 417 4941
rect 383 4839 417 4873
rect 383 4771 417 4805
rect 383 4703 417 4737
rect 383 4635 417 4669
rect 383 4567 417 4601
rect 383 4499 417 4533
rect 383 4431 417 4465
rect 383 4363 417 4397
rect 383 4295 417 4329
rect 383 4227 417 4261
rect 383 4159 417 4193
rect 383 4091 417 4125
rect 383 4023 417 4057
rect 383 3955 417 3989
rect 383 3887 417 3921
rect 383 3819 417 3853
rect 383 3751 417 3785
rect 383 3683 417 3717
rect 383 3615 417 3649
rect 383 3547 417 3581
rect 383 3479 417 3513
rect 383 3411 417 3445
rect 383 3343 417 3377
rect 383 3275 417 3309
rect 383 3207 417 3241
rect 383 3139 417 3173
rect 383 3071 417 3105
rect 383 3003 417 3037
rect 383 2935 417 2969
rect 383 2867 417 2901
rect 383 2799 417 2833
rect 383 2731 417 2765
rect 383 2663 417 2697
rect 383 2595 417 2629
rect 383 2527 417 2561
rect 383 2459 417 2493
rect 383 2391 417 2425
rect 383 2323 417 2357
rect 383 2255 417 2289
rect 383 2187 417 2221
rect 383 2119 417 2153
rect 383 2051 417 2085
rect 383 1983 417 2017
rect 383 1915 417 1949
rect 383 1847 417 1881
rect 383 1779 417 1813
rect 383 1711 417 1745
rect 383 1643 417 1677
rect 383 1575 417 1609
rect 383 1507 417 1541
rect 383 1439 417 1473
rect 383 1371 417 1405
rect 383 1303 417 1337
rect 383 1235 417 1269
rect 383 1167 417 1201
rect 383 1099 417 1133
rect 383 1031 417 1065
rect 383 963 417 997
rect 383 895 417 929
rect 383 827 417 861
rect 383 759 417 793
rect 383 691 417 725
rect 383 623 417 657
rect 383 555 417 589
rect 383 487 417 521
rect 383 419 417 453
rect 383 351 417 385
rect 383 283 417 317
rect 383 215 417 249
rect 383 147 417 181
rect 383 79 417 113
rect 383 11 417 45
rect 383 -57 417 -23
rect 383 -125 417 -91
rect 383 -193 417 -159
rect 383 -261 417 -227
rect 383 -329 417 -295
rect 383 -397 417 -363
rect 22463 5779 22497 5813
rect 22463 5711 22497 5745
rect 22463 5643 22497 5677
rect 22463 5575 22497 5609
rect 22463 5507 22497 5541
rect 22463 5439 22497 5473
rect 22463 5371 22497 5405
rect 22463 5303 22497 5337
rect 22463 5235 22497 5269
rect 22463 5167 22497 5201
rect 22463 5099 22497 5133
rect 22463 5031 22497 5065
rect 22463 4963 22497 4997
rect 22463 4895 22497 4929
rect 22463 4827 22497 4861
rect 22463 4759 22497 4793
rect 22463 4691 22497 4725
rect 22463 4623 22497 4657
rect 22463 4555 22497 4589
rect 22463 4487 22497 4521
rect 22463 4419 22497 4453
rect 22463 4351 22497 4385
rect 22463 4283 22497 4317
rect 22463 4215 22497 4249
rect 22463 4147 22497 4181
rect 22463 4079 22497 4113
rect 22463 4011 22497 4045
rect 22463 3943 22497 3977
rect 22463 3875 22497 3909
rect 22463 3807 22497 3841
rect 22463 3739 22497 3773
rect 22463 3671 22497 3705
rect 22463 3603 22497 3637
rect 22463 3535 22497 3569
rect 22463 3467 22497 3501
rect 22463 3399 22497 3433
rect 22463 3331 22497 3365
rect 22463 3263 22497 3297
rect 22463 3195 22497 3229
rect 22463 3127 22497 3161
rect 22463 3059 22497 3093
rect 22463 2991 22497 3025
rect 22463 2923 22497 2957
rect 22463 2855 22497 2889
rect 22463 2787 22497 2821
rect 22463 2719 22497 2753
rect 22463 2651 22497 2685
rect 22463 2583 22497 2617
rect 22463 2515 22497 2549
rect 22463 2447 22497 2481
rect 22463 2379 22497 2413
rect 22463 2311 22497 2345
rect 22463 2243 22497 2277
rect 22463 2175 22497 2209
rect 22463 2107 22497 2141
rect 22463 2039 22497 2073
rect 22463 1971 22497 2005
rect 22463 1903 22497 1937
rect 22463 1835 22497 1869
rect 22463 1767 22497 1801
rect 22463 1699 22497 1733
rect 22463 1631 22497 1665
rect 22463 1563 22497 1597
rect 22463 1495 22497 1529
rect 22463 1427 22497 1461
rect 22463 1359 22497 1393
rect 22463 1291 22497 1325
rect 22463 1223 22497 1257
rect 22463 1155 22497 1189
rect 22463 1087 22497 1121
rect 22463 1019 22497 1053
rect 22463 951 22497 985
rect 22463 883 22497 917
rect 22463 815 22497 849
rect 22463 747 22497 781
rect 22463 679 22497 713
rect 22463 611 22497 645
rect 22463 543 22497 577
rect 22463 475 22497 509
rect 22463 407 22497 441
rect 22463 339 22497 373
rect 22463 271 22497 305
rect 22463 203 22497 237
rect 22463 135 22497 169
rect 22463 67 22497 101
rect 22463 -1 22497 33
rect 22463 -69 22497 -35
rect 22463 -137 22497 -103
rect 22463 -205 22497 -171
rect 22463 -273 22497 -239
rect 22463 -341 22497 -307
rect 383 -465 417 -431
rect 19140 -423 19240 -374
rect 383 -533 417 -499
rect 383 -601 417 -567
rect 1500 -493 1600 -444
rect 1500 -527 1533 -493
rect 1567 -527 1600 -493
rect 1500 -576 1600 -527
rect 1680 -493 1780 -444
rect 1680 -527 1713 -493
rect 1747 -527 1780 -493
rect 19140 -457 19173 -423
rect 19207 -457 19240 -423
rect 19140 -506 19240 -457
rect 21110 -433 21210 -384
rect 21110 -467 21143 -433
rect 21177 -467 21210 -433
rect 21110 -516 21210 -467
rect 21480 -433 21580 -384
rect 21480 -467 21513 -433
rect 21547 -467 21580 -433
rect 21480 -516 21580 -467
rect 22463 -409 22497 -375
rect 22463 -477 22497 -443
rect 1680 -576 1780 -527
rect 22463 -545 22497 -511
rect 383 -683 417 -635
rect 22463 -613 22497 -579
rect 22463 -683 22497 -647
rect 383 -717 475 -683
rect 509 -717 543 -683
rect 577 -717 611 -683
rect 645 -717 679 -683
rect 713 -717 747 -683
rect 781 -717 815 -683
rect 849 -717 883 -683
rect 917 -717 951 -683
rect 985 -717 1019 -683
rect 1053 -717 1087 -683
rect 1121 -717 1155 -683
rect 1189 -717 1223 -683
rect 1257 -717 1291 -683
rect 1325 -717 1359 -683
rect 1393 -717 1427 -683
rect 1461 -717 1495 -683
rect 1529 -717 1563 -683
rect 1597 -717 1631 -683
rect 1665 -717 1699 -683
rect 1733 -717 1767 -683
rect 1801 -717 1835 -683
rect 1869 -717 1903 -683
rect 1937 -717 1971 -683
rect 2005 -717 2039 -683
rect 2073 -717 2107 -683
rect 2141 -717 2175 -683
rect 2209 -717 2243 -683
rect 2277 -717 2311 -683
rect 2345 -717 2379 -683
rect 2413 -717 2447 -683
rect 2481 -717 2515 -683
rect 2549 -717 2583 -683
rect 2617 -717 2651 -683
rect 2685 -717 2719 -683
rect 2753 -717 2787 -683
rect 2821 -717 2855 -683
rect 2889 -717 2923 -683
rect 2957 -717 2991 -683
rect 3025 -717 3059 -683
rect 3093 -717 3127 -683
rect 3161 -717 3195 -683
rect 3229 -717 3263 -683
rect 3297 -717 3331 -683
rect 3365 -717 3399 -683
rect 3433 -717 3467 -683
rect 3501 -717 3535 -683
rect 3569 -717 3603 -683
rect 3637 -717 3671 -683
rect 3705 -717 3739 -683
rect 3773 -717 3807 -683
rect 3841 -717 3875 -683
rect 3909 -717 3943 -683
rect 3977 -717 4011 -683
rect 4045 -717 4079 -683
rect 4113 -717 4147 -683
rect 4181 -717 4215 -683
rect 4249 -717 4283 -683
rect 4317 -717 4351 -683
rect 4385 -717 4419 -683
rect 4453 -717 4487 -683
rect 4521 -717 4555 -683
rect 4589 -717 4623 -683
rect 4657 -717 4691 -683
rect 4725 -717 4759 -683
rect 4793 -717 4827 -683
rect 4861 -717 4895 -683
rect 4929 -717 4963 -683
rect 4997 -717 5031 -683
rect 5065 -717 5099 -683
rect 5133 -717 5167 -683
rect 5201 -717 5235 -683
rect 5269 -717 5303 -683
rect 5337 -717 5371 -683
rect 5405 -717 5439 -683
rect 5473 -717 5507 -683
rect 5541 -717 5575 -683
rect 5609 -717 5643 -683
rect 5677 -717 5711 -683
rect 5745 -717 5779 -683
rect 5813 -717 5847 -683
rect 5881 -717 5915 -683
rect 5949 -717 5983 -683
rect 6017 -717 6051 -683
rect 6085 -717 6119 -683
rect 6153 -717 6187 -683
rect 6221 -717 6255 -683
rect 6289 -717 6323 -683
rect 6357 -717 6391 -683
rect 6425 -717 6459 -683
rect 6493 -717 6527 -683
rect 6561 -717 6595 -683
rect 6629 -717 6663 -683
rect 6697 -717 6731 -683
rect 6765 -717 6799 -683
rect 6833 -717 6867 -683
rect 6901 -717 6935 -683
rect 6969 -717 7003 -683
rect 7037 -717 7071 -683
rect 7105 -717 7139 -683
rect 7173 -717 7207 -683
rect 7241 -717 7275 -683
rect 7309 -717 7343 -683
rect 7377 -717 7411 -683
rect 7445 -717 7479 -683
rect 7513 -717 7547 -683
rect 7581 -717 7615 -683
rect 7649 -717 7683 -683
rect 7717 -717 7751 -683
rect 7785 -717 7819 -683
rect 7853 -717 7887 -683
rect 7921 -717 7955 -683
rect 7989 -717 8023 -683
rect 8057 -717 8091 -683
rect 8125 -717 8159 -683
rect 8193 -717 8227 -683
rect 8261 -717 8295 -683
rect 8329 -717 8363 -683
rect 8397 -717 8431 -683
rect 8465 -717 8499 -683
rect 8533 -717 8567 -683
rect 8601 -717 8635 -683
rect 8669 -717 8703 -683
rect 8737 -717 8771 -683
rect 8805 -717 8839 -683
rect 8873 -717 8907 -683
rect 8941 -717 8975 -683
rect 9009 -717 9043 -683
rect 9077 -717 9111 -683
rect 9145 -717 9179 -683
rect 9213 -717 9247 -683
rect 9281 -717 9315 -683
rect 9349 -717 9383 -683
rect 9417 -717 9451 -683
rect 9485 -717 9519 -683
rect 9553 -717 9587 -683
rect 9621 -717 9655 -683
rect 9689 -717 9723 -683
rect 9757 -717 9791 -683
rect 9825 -717 9859 -683
rect 9893 -717 9927 -683
rect 9961 -717 9995 -683
rect 10029 -717 10063 -683
rect 10097 -717 10131 -683
rect 10165 -717 10199 -683
rect 10233 -717 10267 -683
rect 10301 -717 10335 -683
rect 10369 -717 10403 -683
rect 10437 -717 10471 -683
rect 10505 -717 10539 -683
rect 10573 -717 10607 -683
rect 10641 -717 10675 -683
rect 10709 -717 10743 -683
rect 10777 -717 10811 -683
rect 10845 -717 10879 -683
rect 10913 -717 10947 -683
rect 10981 -717 11015 -683
rect 11049 -717 11083 -683
rect 11117 -717 11151 -683
rect 11185 -717 11219 -683
rect 11253 -717 11287 -683
rect 11321 -717 11355 -683
rect 11389 -717 11423 -683
rect 11457 -717 11491 -683
rect 11525 -717 11559 -683
rect 11593 -717 11627 -683
rect 11661 -717 11695 -683
rect 11729 -717 11763 -683
rect 11797 -717 11831 -683
rect 11865 -717 11899 -683
rect 11933 -717 11967 -683
rect 12001 -717 12035 -683
rect 12069 -717 12103 -683
rect 12137 -717 12171 -683
rect 12205 -717 12239 -683
rect 12273 -717 12307 -683
rect 12341 -717 12375 -683
rect 12409 -717 12443 -683
rect 12477 -717 12511 -683
rect 12545 -717 12579 -683
rect 12613 -717 12647 -683
rect 12681 -717 12715 -683
rect 12749 -717 12783 -683
rect 12817 -717 12851 -683
rect 12885 -717 12919 -683
rect 12953 -717 12987 -683
rect 13021 -717 13055 -683
rect 13089 -717 13123 -683
rect 13157 -717 13191 -683
rect 13225 -717 13259 -683
rect 13293 -717 13327 -683
rect 13361 -717 13395 -683
rect 13429 -717 13463 -683
rect 13497 -717 13531 -683
rect 13565 -717 13599 -683
rect 13633 -717 13667 -683
rect 13701 -717 13735 -683
rect 13769 -717 13803 -683
rect 13837 -717 13871 -683
rect 13905 -717 13939 -683
rect 13973 -717 14007 -683
rect 14041 -717 14075 -683
rect 14109 -717 14143 -683
rect 14177 -717 14211 -683
rect 14245 -717 14279 -683
rect 14313 -717 14347 -683
rect 14381 -717 14415 -683
rect 14449 -717 14483 -683
rect 14517 -717 14551 -683
rect 14585 -717 14619 -683
rect 14653 -717 14687 -683
rect 14721 -717 14755 -683
rect 14789 -717 14823 -683
rect 14857 -717 14891 -683
rect 14925 -717 14959 -683
rect 14993 -717 15027 -683
rect 15061 -717 15095 -683
rect 15129 -717 15163 -683
rect 15197 -717 15231 -683
rect 15265 -717 15299 -683
rect 15333 -717 15367 -683
rect 15401 -717 15435 -683
rect 15469 -717 15503 -683
rect 15537 -717 15571 -683
rect 15605 -717 15639 -683
rect 15673 -717 15707 -683
rect 15741 -717 15775 -683
rect 15809 -717 15843 -683
rect 15877 -717 15911 -683
rect 15945 -717 15979 -683
rect 16013 -717 16047 -683
rect 16081 -717 16115 -683
rect 16149 -717 16183 -683
rect 16217 -717 16251 -683
rect 16285 -717 16319 -683
rect 16353 -717 16387 -683
rect 16421 -717 16455 -683
rect 16489 -717 16523 -683
rect 16557 -717 16591 -683
rect 16625 -717 16659 -683
rect 16693 -717 16727 -683
rect 16761 -717 16795 -683
rect 16829 -717 16863 -683
rect 16897 -717 16931 -683
rect 16965 -717 16999 -683
rect 17033 -717 17067 -683
rect 17101 -717 17135 -683
rect 17169 -717 17203 -683
rect 17237 -717 17271 -683
rect 17305 -717 17339 -683
rect 17373 -717 17407 -683
rect 17441 -717 17475 -683
rect 17509 -717 17543 -683
rect 17577 -717 17611 -683
rect 17645 -717 17679 -683
rect 17713 -717 17747 -683
rect 17781 -717 17815 -683
rect 17849 -717 17883 -683
rect 17917 -717 17951 -683
rect 17985 -717 18019 -683
rect 18053 -717 18087 -683
rect 18121 -717 18155 -683
rect 18189 -717 18223 -683
rect 18257 -717 18291 -683
rect 18325 -717 18359 -683
rect 18393 -717 18427 -683
rect 18461 -717 18495 -683
rect 18529 -717 18563 -683
rect 18597 -717 18631 -683
rect 18665 -717 18699 -683
rect 18733 -717 18767 -683
rect 18801 -717 18835 -683
rect 18869 -717 18903 -683
rect 18937 -717 18971 -683
rect 19005 -717 19039 -683
rect 19073 -717 19107 -683
rect 19141 -717 19175 -683
rect 19209 -717 19243 -683
rect 19277 -717 19311 -683
rect 19345 -717 19379 -683
rect 19413 -717 19447 -683
rect 19481 -717 19515 -683
rect 19549 -717 19583 -683
rect 19617 -717 19651 -683
rect 19685 -717 19719 -683
rect 19753 -717 19787 -683
rect 19821 -717 19855 -683
rect 19889 -717 19923 -683
rect 19957 -717 19991 -683
rect 20025 -717 20059 -683
rect 20093 -717 20127 -683
rect 20161 -717 20195 -683
rect 20229 -717 20263 -683
rect 20297 -717 20331 -683
rect 20365 -717 20399 -683
rect 20433 -717 20467 -683
rect 20501 -717 20535 -683
rect 20569 -717 20603 -683
rect 20637 -717 20671 -683
rect 20705 -717 20739 -683
rect 20773 -717 20807 -683
rect 20841 -717 20875 -683
rect 20909 -717 20943 -683
rect 20977 -717 21011 -683
rect 21045 -717 21079 -683
rect 21113 -717 21147 -683
rect 21181 -717 21215 -683
rect 21249 -717 21283 -683
rect 21317 -717 21351 -683
rect 21385 -717 21419 -683
rect 21453 -717 21487 -683
rect 21521 -717 21555 -683
rect 21589 -717 21623 -683
rect 21657 -717 21691 -683
rect 21725 -717 21759 -683
rect 21793 -717 21827 -683
rect 21861 -717 21895 -683
rect 21929 -717 21963 -683
rect 21997 -717 22031 -683
rect 22065 -717 22099 -683
rect 22133 -717 22167 -683
rect 22201 -717 22235 -683
rect 22269 -717 22303 -683
rect 22337 -717 22371 -683
rect 22405 -717 22497 -683
<< viali >>
rect 1030 21408 1064 21442
rect 1102 21408 1109 21442
rect 1109 21408 1136 21442
rect 1174 21408 1177 21442
rect 1177 21408 1208 21442
rect 1246 21408 1280 21442
rect 7020 21403 7054 21437
rect 7092 21403 7123 21437
rect 7123 21403 7126 21437
rect 7164 21403 7191 21437
rect 7191 21403 7198 21437
rect 7236 21403 7270 21437
rect 2723 12313 2757 12347
rect 2903 12313 2937 12347
rect 5623 12303 5657 12337
rect 5803 12303 5837 12337
rect 14323 10373 14357 10407
rect 1623 5843 1657 5877
rect 19173 -457 19207 -423
rect 21143 -467 21177 -433
<< metal1 >>
rect 1010 21442 1310 21860
rect 1010 21408 1030 21442
rect 1064 21408 1102 21442
rect 1136 21408 1174 21442
rect 1208 21408 1246 21442
rect 1280 21408 1310 21442
rect 1010 20970 1310 21408
rect 1890 20920 2190 21860
rect 2800 20920 3100 21860
rect 3680 20910 3980 21860
rect 4590 20910 4890 21860
rect 5490 20940 5790 21860
rect 6390 20920 6690 21860
rect 7000 21437 7300 21860
rect 7000 21403 7020 21437
rect 7054 21403 7092 21437
rect 7126 21403 7164 21437
rect 7198 21403 7236 21437
rect 7270 21403 7300 21437
rect 7000 20910 7300 21403
rect 8190 21320 8490 21860
rect 8970 21280 9270 21340
rect 9790 21270 10090 21860
rect 10580 21270 10880 21340
rect 11360 21310 11660 21860
rect 7460 18030 8210 18190
rect 7460 17670 7510 18030
rect 8060 17940 8210 18030
rect 8060 17670 8490 17940
rect 9240 17930 10900 17950
rect 12080 17930 12460 18240
rect 10560 17670 10850 17930
rect 8190 17650 8490 17670
rect 9240 17650 10850 17670
rect 10830 17630 10850 17650
rect 10800 17400 10850 17630
rect 12460 17310 12600 17620
rect 7490 15880 8060 16090
rect 930 12740 1290 13120
rect 2650 12740 3010 13120
rect 4090 12740 4450 13120
rect 5550 12740 5910 13120
rect 7390 12740 7750 13120
rect 10860 12606 11010 12640
rect 10860 12554 10874 12606
rect 10926 12554 10954 12606
rect 11006 12554 11010 12606
rect 10860 12520 11010 12554
rect 930 12060 1290 12460
rect 2650 12347 3010 12460
rect 2650 12313 2723 12347
rect 2757 12313 2903 12347
rect 2937 12313 3010 12347
rect 2650 12060 3010 12313
rect 4090 12050 4450 12460
rect 5550 12337 5910 12460
rect 5550 12303 5623 12337
rect 5657 12303 5803 12337
rect 5837 12303 5910 12337
rect 5550 12050 5910 12303
rect 7390 12060 7750 12460
rect 9330 11580 9950 11620
rect 10890 10770 11010 12520
rect 10890 10736 11090 10770
rect 10890 10684 10909 10736
rect 10961 10684 11019 10736
rect 11071 10684 11090 10736
rect 10890 10650 11090 10684
rect 14190 10407 14490 10460
rect 14190 10373 14323 10407
rect 14357 10373 14490 10407
rect 10490 10110 11890 10270
rect 11710 9650 11890 10110
rect 11710 9640 12120 9650
rect 11350 9580 12120 9640
rect 14190 9630 14490 10373
rect 15300 9640 15610 10460
rect 16370 9640 16680 10460
rect 18870 9710 19170 9760
rect 19720 9710 20020 10450
rect 20560 9710 20860 10290
rect 21400 9710 21700 10430
rect 15300 9630 15600 9640
rect 16370 9630 16670 9640
rect 17200 9630 17510 9640
rect 960 6380 1260 6750
rect 1570 6380 1870 6750
rect 2730 6380 3030 6750
rect 3890 6380 4190 6750
rect 5050 6380 5350 6750
rect 6210 6380 6510 6750
rect 7380 6380 7680 6750
rect 1570 5877 1870 6070
rect 1570 5843 1623 5877
rect 1657 5843 1870 5877
rect 1570 5250 1870 5843
rect 2720 5260 3020 6080
rect 18930 220 19230 260
rect 19710 220 20010 260
rect 20550 220 20850 260
rect 21470 220 21770 260
rect 3160 30 3520 40
rect 1430 20 1730 30
rect 1430 10 1790 20
rect 2250 10 2550 30
rect 3160 10 3590 30
rect 4350 10 4650 30
rect 5220 10 5670 30
rect 6530 10 6830 40
rect 1430 0 6830 10
rect 1430 -680 1790 0
rect 3160 -720 3520 0
rect 5220 -730 5580 0
rect 8860 -370 9170 -320
rect 11130 -370 11340 -290
rect 8860 -720 9220 -370
rect 10980 -720 11340 -370
rect 14710 -370 14850 -290
rect 17070 -360 17270 -290
rect 14710 -720 15070 -370
rect 17070 -720 17430 -360
rect 19080 -423 19440 220
rect 19080 -457 19173 -423
rect 19207 -457 19440 -423
rect 19080 -720 19440 -457
rect 21040 -433 21400 220
rect 21040 -467 21143 -433
rect 21177 -467 21400 -433
rect 21040 -920 21400 -467
<< via1 >>
rect 10874 12554 10926 12606
rect 10954 12554 11006 12606
rect 10909 10684 10961 10736
rect 11019 10684 11071 10736
<< metal2 >>
rect 8180 12608 11010 12640
rect 8180 12552 8197 12608
rect 8253 12552 8307 12608
rect 8363 12606 11010 12608
rect 8363 12554 10874 12606
rect 10926 12554 10954 12606
rect 11006 12554 11010 12606
rect 8363 12552 11010 12554
rect 8180 12520 11010 12552
rect 8440 11328 8560 11350
rect 8440 11272 8472 11328
rect 8528 11310 8560 11328
rect 8528 11280 8830 11310
rect 8528 11272 9890 11280
rect 8440 11250 9890 11272
rect 8770 11220 9890 11250
rect 8640 11190 8740 11210
rect 8640 11188 8860 11190
rect 8640 11132 8662 11188
rect 8718 11132 8860 11188
rect 8640 11130 8860 11132
rect 8640 11110 8740 11130
rect 21290 10770 21370 11480
rect 10890 10738 11090 10770
rect 10890 10682 10907 10738
rect 10963 10682 11017 10738
rect 11073 10682 11090 10738
rect 10890 10650 11090 10682
rect 21170 10738 21370 10770
rect 21170 10682 21187 10738
rect 21243 10682 21297 10738
rect 21353 10682 21370 10738
rect 21170 10650 21370 10682
rect 8270 9278 8350 9290
rect 8270 9222 8282 9278
rect 8338 9222 8350 9278
rect 8270 9210 8350 9222
<< via2 >>
rect 8197 12552 8253 12608
rect 8307 12552 8363 12608
rect 8472 11272 8528 11328
rect 8662 11132 8718 11188
rect 10907 10736 10963 10738
rect 10907 10684 10909 10736
rect 10909 10684 10961 10736
rect 10961 10684 10963 10736
rect 10907 10682 10963 10684
rect 11017 10736 11073 10738
rect 11017 10684 11019 10736
rect 11019 10684 11071 10736
rect 11071 10684 11073 10736
rect 11017 10682 11073 10684
rect 21187 10682 21243 10738
rect 21297 10682 21353 10738
rect 8282 9222 8338 9278
<< metal3 >>
rect -60 21782 80 21820
rect -60 21718 -22 21782
rect 42 21718 80 21782
rect -60 15242 80 21718
rect 7650 21782 7770 21790
rect 7650 21718 7678 21782
rect 7742 21718 7770 21782
rect 220 21583 360 21626
rect 220 21519 258 21583
rect 322 21519 360 21583
rect 220 15422 360 21519
rect 7410 21582 7530 21620
rect 7410 21518 7438 21582
rect 7502 21518 7530 21582
rect 7410 21360 7530 21518
rect 7650 21360 7770 21718
rect 8040 21777 8160 21790
rect 8040 21713 8063 21777
rect 8127 21713 8160 21777
rect 7840 21582 7960 21620
rect 7840 21518 7868 21582
rect 7932 21518 7960 21582
rect 7840 21240 7960 21518
rect 8040 21240 8160 21713
rect 450 21127 570 21160
rect 450 21063 478 21127
rect 542 21063 570 21127
rect 450 15602 570 21063
rect 10960 16012 11080 16980
rect 10960 15948 10988 16012
rect 11052 15948 11080 16012
rect 10960 15920 11080 15948
rect 11430 16012 11550 16040
rect 11430 15948 11458 16012
rect 11522 15948 11550 16012
rect 10960 15772 11080 15800
rect 10960 15708 10988 15772
rect 11052 15708 11080 15772
rect 10960 15680 11080 15708
rect 11250 15772 11370 15800
rect 11250 15708 11278 15772
rect 11342 15708 11370 15772
rect 450 15538 478 15602
rect 542 15538 570 15602
rect 450 15510 570 15538
rect 3450 15597 3590 15630
rect 3450 15533 3493 15597
rect 3557 15533 3590 15597
rect 220 15358 258 15422
rect 322 15358 360 15422
rect 220 15330 360 15358
rect 3250 15422 3390 15450
rect 3250 15358 3288 15422
rect 3352 15358 3390 15422
rect -60 15178 -22 15242
rect 42 15178 80 15242
rect -60 15150 80 15178
rect 1460 15242 1600 15260
rect 1460 15178 1498 15242
rect 1562 15178 1600 15242
rect 1460 12150 1600 15178
rect 3250 12410 3390 15358
rect 3450 13322 3590 15533
rect 7390 14122 7510 15640
rect 7630 14387 7750 15590
rect 7630 14323 7658 14387
rect 7722 14323 7750 14387
rect 7630 14277 7750 14323
rect 7630 14213 7658 14277
rect 7722 14213 7750 14277
rect 7630 14190 7750 14213
rect 10590 14287 10830 14310
rect 10590 14223 10618 14287
rect 10682 14223 10738 14287
rect 10802 14223 10830 14287
rect 10590 14190 10830 14223
rect 10950 14282 11190 14310
rect 10950 14218 10978 14282
rect 11042 14218 11098 14282
rect 11162 14218 11190 14282
rect 10950 14190 11190 14218
rect 7390 14058 7418 14122
rect 7482 14058 7510 14122
rect 7390 14002 7510 14058
rect 7390 13938 7418 14002
rect 7482 13938 7510 14002
rect 7390 13910 7510 13938
rect 10410 14002 10650 14030
rect 10410 13938 10438 14002
rect 10502 13938 10558 14002
rect 10622 13938 10650 14002
rect 10410 13910 10650 13938
rect 3450 13258 3488 13322
rect 3552 13258 3590 13322
rect 3450 13230 3590 13258
rect 8440 13322 8560 13350
rect 8440 13258 8468 13322
rect 8532 13258 8560 13322
rect 8180 12612 8380 12640
rect 8180 12548 8193 12612
rect 8257 12548 8303 12612
rect 8367 12548 8380 12612
rect 8180 12520 8380 12548
rect 3240 12280 3400 12410
rect 3250 12150 3390 12280
rect 8260 12243 8380 12280
rect 8260 12179 8288 12243
rect 8352 12179 8380 12243
rect 8260 10199 8380 12179
rect 8440 11328 8560 13258
rect 8440 11272 8472 11328
rect 8528 11272 8560 11328
rect 8440 11250 8560 11272
rect 8630 12432 8750 12460
rect 8630 12368 8658 12432
rect 8722 12368 8750 12432
rect 8630 11188 8750 12368
rect 8630 11132 8662 11188
rect 8718 11132 8750 11188
rect 8630 11110 8750 11132
rect 10530 10382 10650 13910
rect 10710 10562 10830 14190
rect 10890 14002 11010 14030
rect 10890 13938 10918 14002
rect 10982 13938 11010 14002
rect 10890 10932 11010 13938
rect 11070 11132 11190 14190
rect 11250 11312 11370 15708
rect 11430 11492 11550 15948
rect 12280 15772 12400 21200
rect 12280 15708 12308 15772
rect 12372 15708 12400 15772
rect 12280 15680 12400 15708
rect 12530 14200 12630 14300
rect 11430 11428 11458 11492
rect 11522 11428 11550 11492
rect 11430 11400 11550 11428
rect 18760 11492 18880 11520
rect 18760 11428 18788 11492
rect 18852 11428 18880 11492
rect 11250 11248 11278 11312
rect 11342 11248 11370 11312
rect 11250 11220 11370 11248
rect 18520 11312 18640 11340
rect 18520 11248 18548 11312
rect 18612 11248 18640 11312
rect 11070 11068 11098 11132
rect 11162 11068 11190 11132
rect 11070 11040 11190 11068
rect 18140 11132 18260 11160
rect 18140 11068 18168 11132
rect 18232 11068 18260 11132
rect 10890 10868 10918 10932
rect 10982 10868 11010 10932
rect 10890 10840 11010 10868
rect 17960 10932 18080 10960
rect 17960 10868 17988 10932
rect 18052 10868 18080 10932
rect 10890 10742 11090 10770
rect 10890 10678 10903 10742
rect 10967 10678 11013 10742
rect 11077 10678 11090 10742
rect 10890 10650 11090 10678
rect 10710 10498 10738 10562
rect 10802 10498 10830 10562
rect 10710 10470 10830 10498
rect 13310 10562 13430 10590
rect 13310 10498 13338 10562
rect 13402 10498 13430 10562
rect 10530 10318 10558 10382
rect 10622 10318 10650 10382
rect 10530 10290 10650 10318
rect 13090 10382 13170 10400
rect 13090 10318 13098 10382
rect 13162 10318 13170 10382
rect 13310 10360 13430 10498
rect 13090 10300 13170 10318
rect 8255 10172 8385 10199
rect 8255 10108 8288 10172
rect 8352 10108 8385 10172
rect 8255 10081 8385 10108
rect 8260 10080 8380 10081
rect 450 9552 530 9560
rect 450 9488 458 9552
rect 522 9488 530 9552
rect 450 9480 530 9488
rect 8260 9278 8360 9300
rect 450 9262 530 9270
rect 450 9198 458 9262
rect 522 9198 530 9262
rect 450 9190 530 9198
rect 8260 9222 8282 9278
rect 8338 9222 8360 9278
rect 8260 7110 8360 9222
rect 7460 5410 7950 5510
rect 7460 5210 7790 5310
rect 7690 652 7790 5210
rect 7850 2842 7950 5410
rect 17960 5010 18080 10868
rect 18140 7160 18260 11068
rect 18520 9900 18640 11248
rect 18760 10932 18880 11428
rect 18760 10868 18788 10932
rect 18852 10868 18880 10932
rect 18760 10840 18880 10868
rect 21960 10932 22080 10960
rect 21960 10868 21988 10932
rect 22052 10868 22080 10932
rect 21170 10742 21370 10770
rect 21170 10678 21183 10742
rect 21247 10678 21293 10742
rect 21357 10678 21370 10742
rect 21170 10650 21370 10678
rect 21960 9900 22080 10868
rect 17960 4890 18260 5010
rect 7850 2778 7868 2842
rect 7932 2778 7950 2842
rect 7850 2760 7950 2778
rect 8270 2842 8350 2850
rect 8270 2778 8278 2842
rect 8342 2778 8350 2842
rect 8270 2770 8350 2778
rect 7690 588 7708 652
rect 7772 588 7790 652
rect 7690 570 7790 588
rect 8100 652 8200 670
rect 8100 588 8118 652
rect 8182 588 8200 652
rect 7460 492 7560 510
rect 7460 428 7478 492
rect 7542 428 7560 492
rect 7460 410 7560 428
rect 7940 492 8040 510
rect 7940 428 7958 492
rect 8022 428 8040 492
rect 7460 292 7560 310
rect 7460 228 7478 292
rect 7542 228 7560 292
rect 7460 210 7560 228
rect 7780 292 7880 310
rect 7780 228 7798 292
rect 7862 228 7880 292
rect 7460 -10 7720 90
rect 7460 -578 7560 -100
rect 7620 -418 7720 -10
rect 7780 -219 7880 228
rect 7940 -18 8040 428
rect 8100 200 8200 588
rect 8100 100 8360 200
rect 7940 -82 7958 -18
rect 8022 -82 8040 -18
rect 7940 -100 8040 -82
rect 8270 -18 8350 -10
rect 8270 -82 8278 -18
rect 8342 -82 8350 -18
rect 8270 -90 8350 -82
rect 7780 -283 7798 -219
rect 7862 -283 7880 -219
rect 7780 -306 7880 -283
rect 8261 -219 8359 -196
rect 8261 -283 8278 -219
rect 8342 -283 8359 -219
rect 8261 -306 8359 -283
rect 7620 -482 7638 -418
rect 7702 -482 7720 -418
rect 7620 -500 7720 -482
rect 18380 -418 18480 -90
rect 18380 -482 18398 -418
rect 18462 -482 18480 -418
rect 18380 -500 18480 -482
rect 7460 -642 7478 -578
rect 7542 -642 7560 -578
rect 7460 -660 7560 -642
rect 18680 -578 18780 -90
rect 18680 -642 18698 -578
rect 18762 -642 18780 -578
rect 18680 -660 18780 -642
rect 22340 -1148 22460 2740
rect 22340 -1212 22368 -1148
rect 22432 -1212 22460 -1148
rect 22340 -1230 22460 -1212
<< via3 >>
rect -22 21718 42 21782
rect 7678 21718 7742 21782
rect 258 21519 322 21583
rect 7438 21518 7502 21582
rect 8063 21713 8127 21777
rect 7868 21518 7932 21582
rect 478 21063 542 21127
rect 10988 15948 11052 16012
rect 11458 15948 11522 16012
rect 10988 15708 11052 15772
rect 11278 15708 11342 15772
rect 478 15538 542 15602
rect 3493 15533 3557 15597
rect 258 15358 322 15422
rect 3288 15358 3352 15422
rect -22 15178 42 15242
rect 1498 15178 1562 15242
rect 7658 14323 7722 14387
rect 7658 14213 7722 14277
rect 10618 14223 10682 14287
rect 10738 14223 10802 14287
rect 10978 14218 11042 14282
rect 11098 14218 11162 14282
rect 7418 14058 7482 14122
rect 7418 13938 7482 14002
rect 10438 13938 10502 14002
rect 10558 13938 10622 14002
rect 3488 13258 3552 13322
rect 8468 13258 8532 13322
rect 8193 12608 8257 12612
rect 8193 12552 8197 12608
rect 8197 12552 8253 12608
rect 8253 12552 8257 12608
rect 8193 12548 8257 12552
rect 8303 12608 8367 12612
rect 8303 12552 8307 12608
rect 8307 12552 8363 12608
rect 8363 12552 8367 12608
rect 8303 12548 8367 12552
rect 8288 12179 8352 12243
rect 8658 12368 8722 12432
rect 10918 13938 10982 14002
rect 12308 15708 12372 15772
rect 11458 11428 11522 11492
rect 18788 11428 18852 11492
rect 11278 11248 11342 11312
rect 18548 11248 18612 11312
rect 11098 11068 11162 11132
rect 18168 11068 18232 11132
rect 10918 10868 10982 10932
rect 17988 10868 18052 10932
rect 10903 10738 10967 10742
rect 10903 10682 10907 10738
rect 10907 10682 10963 10738
rect 10963 10682 10967 10738
rect 10903 10678 10967 10682
rect 11013 10738 11077 10742
rect 11013 10682 11017 10738
rect 11017 10682 11073 10738
rect 11073 10682 11077 10738
rect 11013 10678 11077 10682
rect 10738 10498 10802 10562
rect 13338 10498 13402 10562
rect 10558 10318 10622 10382
rect 13098 10318 13162 10382
rect 8288 10108 8352 10172
rect 458 9488 522 9552
rect 458 9198 522 9262
rect 18788 10868 18852 10932
rect 21988 10868 22052 10932
rect 21183 10738 21247 10742
rect 21183 10682 21187 10738
rect 21187 10682 21243 10738
rect 21243 10682 21247 10738
rect 21183 10678 21247 10682
rect 21293 10738 21357 10742
rect 21293 10682 21297 10738
rect 21297 10682 21353 10738
rect 21353 10682 21357 10738
rect 21293 10678 21357 10682
rect 7868 2778 7932 2842
rect 8278 2778 8342 2842
rect 7708 588 7772 652
rect 8118 588 8182 652
rect 7478 428 7542 492
rect 7958 428 8022 492
rect 7478 228 7542 292
rect 7798 228 7862 292
rect 7958 -82 8022 -18
rect 8278 -82 8342 -18
rect 7798 -283 7862 -219
rect 8278 -283 8342 -219
rect 7638 -482 7702 -418
rect 18398 -482 18462 -418
rect 7478 -642 7542 -578
rect 18698 -642 18762 -578
rect 22368 -1212 22432 -1148
<< metal4 >>
rect -60 21782 8160 21810
rect -60 21718 -22 21782
rect 42 21718 7678 21782
rect 7742 21777 8160 21782
rect 7742 21718 8063 21777
rect -60 21713 8063 21718
rect 8127 21713 8160 21777
rect -60 21681 8160 21713
rect -60 21680 80 21681
rect 219 21583 7960 21621
rect 219 21519 258 21583
rect 322 21582 7960 21583
rect 322 21519 7438 21582
rect 219 21518 7438 21519
rect 7502 21518 7868 21582
rect 7932 21518 7960 21582
rect 219 21481 7960 21518
rect 450 21127 570 21230
rect 450 21063 478 21127
rect 542 21063 570 21127
rect 450 21030 570 21063
rect 10960 16012 11550 16040
rect 10960 15948 10988 16012
rect 11052 15948 11458 16012
rect 11522 15948 11550 16012
rect 10960 15920 11550 15948
rect 10960 15772 12400 15800
rect 10960 15708 10988 15772
rect 11052 15708 11278 15772
rect 11342 15708 12308 15772
rect 12372 15708 12400 15772
rect 10960 15680 12400 15708
rect 450 15602 3590 15630
rect 450 15538 478 15602
rect 542 15597 3590 15602
rect 542 15538 3493 15597
rect 450 15533 3493 15538
rect 3557 15533 3590 15597
rect 450 15510 3590 15533
rect 220 15422 3390 15450
rect 220 15358 258 15422
rect 322 15358 3288 15422
rect 3352 15358 3390 15422
rect 220 15330 3390 15358
rect -60 15242 1600 15270
rect -60 15178 -22 15242
rect 42 15178 1498 15242
rect 1562 15178 1600 15242
rect -60 15150 1600 15178
rect 7630 14387 7750 14410
rect 7630 14323 7658 14387
rect 7722 14370 7750 14387
rect 7722 14323 12650 14370
rect 7630 14287 12650 14323
rect 7630 14277 10618 14287
rect 7630 14213 7658 14277
rect 7722 14223 10618 14277
rect 10682 14223 10738 14287
rect 10802 14282 12650 14287
rect 10802 14223 10978 14282
rect 7722 14218 10978 14223
rect 11042 14218 11098 14282
rect 11162 14218 12650 14282
rect 7722 14213 12650 14218
rect 7630 14190 12650 14213
rect 7390 14122 7510 14150
rect 7390 14058 7418 14122
rect 7482 14090 7510 14122
rect 7482 14058 12830 14090
rect 7390 14002 12830 14058
rect 7390 13938 7418 14002
rect 7482 13938 10438 14002
rect 10502 13938 10558 14002
rect 10622 13938 10918 14002
rect 10982 13938 12830 14002
rect 7390 13910 12830 13938
rect 3450 13322 8560 13350
rect 3450 13258 3488 13322
rect 3552 13258 8468 13322
rect 8532 13258 8560 13322
rect 3450 13230 8560 13258
rect 250 12612 8380 12640
rect 250 12548 8193 12612
rect 8257 12548 8303 12612
rect 8367 12548 8380 12612
rect 250 12520 8380 12548
rect 250 12432 8750 12460
rect 250 12368 8658 12432
rect 8722 12368 8750 12432
rect 250 12340 8750 12368
rect 290 12270 8381 12271
rect 250 12243 8381 12270
rect 250 12179 8288 12243
rect 8352 12179 8381 12243
rect 250 12151 8381 12179
rect 250 12150 350 12151
rect 11430 11492 18880 11520
rect 11430 11428 11458 11492
rect 11522 11428 18788 11492
rect 18852 11428 18880 11492
rect 11430 11400 18880 11428
rect 11250 11312 18640 11340
rect 11250 11248 11278 11312
rect 11342 11248 18548 11312
rect 18612 11248 18640 11312
rect 11250 11220 18640 11248
rect 11070 11132 18260 11160
rect 11070 11068 11098 11132
rect 11162 11068 18168 11132
rect 18232 11068 18260 11132
rect 11070 11040 18260 11068
rect 10890 10932 18080 10960
rect 10890 10868 10918 10932
rect 10982 10868 17988 10932
rect 18052 10868 18080 10932
rect 10890 10840 18080 10868
rect 18760 10932 22080 10960
rect 18760 10868 18788 10932
rect 18852 10868 21988 10932
rect 22052 10868 22080 10932
rect 18760 10840 22080 10868
rect 10890 10742 21370 10770
rect 10890 10678 10903 10742
rect 10967 10678 11013 10742
rect 11077 10678 21183 10742
rect 21247 10678 21293 10742
rect 21357 10678 21370 10742
rect 10890 10650 21370 10678
rect 10710 10562 13430 10590
rect 10710 10498 10738 10562
rect 10802 10498 13338 10562
rect 13402 10498 13430 10562
rect 10710 10470 13430 10498
rect 10530 10382 13180 10410
rect 10530 10318 10558 10382
rect 10622 10318 13098 10382
rect 13162 10318 13180 10382
rect 10530 10290 13180 10318
rect 8260 10172 8380 10200
rect 8260 10108 8288 10172
rect 8352 10108 8380 10172
rect 8260 10080 8380 10108
rect 230 9552 540 9570
rect 230 9488 458 9552
rect 522 9488 540 9552
rect 230 9470 540 9488
rect 230 9262 540 9280
rect 230 9198 458 9262
rect 522 9198 540 9262
rect 230 9180 540 9198
rect 430 5500 780 5600
rect 7850 2842 8360 2860
rect 7850 2778 7868 2842
rect 7932 2778 8278 2842
rect 8342 2778 8360 2842
rect 7850 2760 8360 2778
rect 7690 652 8200 670
rect 7690 588 7708 652
rect 7772 588 8118 652
rect 8182 588 8200 652
rect 7690 570 8200 588
rect 7460 492 8040 510
rect 7460 428 7478 492
rect 7542 428 7958 492
rect 8022 428 8040 492
rect 7460 410 8040 428
rect 7460 292 7880 310
rect 7460 228 7478 292
rect 7542 228 7798 292
rect 7862 228 7880 292
rect 7460 210 7880 228
rect 7940 -18 8360 0
rect 7940 -82 7958 -18
rect 8022 -82 8278 -18
rect 8342 -82 8360 -18
rect 7940 -100 8360 -82
rect 7779 -219 8360 -201
rect 7779 -283 7798 -219
rect 7862 -283 8278 -219
rect 8342 -283 8360 -219
rect 7779 -301 8360 -283
rect 7620 -418 18480 -400
rect 7620 -482 7638 -418
rect 7702 -482 18398 -418
rect 18462 -482 18480 -418
rect 7620 -500 18480 -482
rect 7460 -578 18780 -560
rect 7460 -642 7478 -578
rect 7542 -642 18698 -578
rect 18762 -642 18780 -578
rect 7460 -660 18780 -642
rect 22340 -1148 22460 -1130
rect 22340 -1212 22368 -1148
rect 22432 -1212 22460 -1148
rect 22340 -1230 22460 -1212
use diff_in_03  diff_in_03_0
timestamp 1757161594
transform 1 0 1450 0 1 7130
box -1010 -673 6910 5260
use diff_in_04  diff_in_04_0
timestamp 1757161594
transform 1 0 18670 0 1 500
box -510 -690 3790 9510
use nmos_08  nmos_08_0
timestamp 1757161594
transform 1 0 8860 0 1 10440
box 0 -26 1634 1212
use nmos_cl_02  nmos_cl_02_1
timestamp 1757161594
transform 1 0 8850 0 1 4950
box -590 -5320 9003 5510
use nmos_cload_01  nmos_cload_01_1
timestamp 1757161594
transform 1 0 1430 0 1 2670
box -770 -2923 6130 3053
use pmos_05  pmos_05_0
timestamp 1757161594
transform 1 0 953 0 1 16170
box -493 -690 6897 5358
use pmos_06  pmos_06_0
timestamp 1757161594
transform 1 0 8130 0 1 18320
box -290 -530 4270 3030
use pmos_07  pmos_07_0
timestamp 1757161594
transform 0 -1 10510 1 0 15280
box -80 -570 2530 2710
<< labels >>
flabel metal4 s 250 12340 350 12440 0 FreeSans 392 0 0 0 Vbias3
port 1 nsew
flabel metal4 s 250 12150 350 12250 0 FreeSans 392 0 0 0 Vbias2
port 2 nsew
<< end >>
