magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -1380 -2320 3380 80
<< nsubdiff >>
rect -1340 17 3340 40
rect -1340 -17 -1227 17
rect -1193 -17 -1159 17
rect -1125 -17 -1091 17
rect -1057 -17 -1023 17
rect -989 -17 -955 17
rect -921 -17 -887 17
rect -853 -17 -819 17
rect -785 -17 -751 17
rect -717 -17 -683 17
rect -649 -17 -615 17
rect -581 -17 -547 17
rect -513 -17 -479 17
rect -445 -17 -411 17
rect -377 -17 -343 17
rect -309 -17 -275 17
rect -241 -17 -207 17
rect -173 -17 -139 17
rect -105 -17 -71 17
rect -37 -17 -3 17
rect 31 -17 65 17
rect 99 -17 133 17
rect 167 -17 201 17
rect 235 -17 269 17
rect 303 -17 337 17
rect 371 -17 405 17
rect 439 -17 473 17
rect 507 -17 541 17
rect 575 -17 609 17
rect 643 -17 677 17
rect 711 -17 745 17
rect 779 -17 813 17
rect 847 -17 881 17
rect 915 -17 949 17
rect 983 -17 1017 17
rect 1051 -17 1085 17
rect 1119 -17 1153 17
rect 1187 -17 1221 17
rect 1255 -17 1289 17
rect 1323 -17 1357 17
rect 1391 -17 1425 17
rect 1459 -17 1493 17
rect 1527 -17 1561 17
rect 1595 -17 1629 17
rect 1663 -17 1697 17
rect 1731 -17 1765 17
rect 1799 -17 1833 17
rect 1867 -17 1901 17
rect 1935 -17 1969 17
rect 2003 -17 2037 17
rect 2071 -17 2105 17
rect 2139 -17 2173 17
rect 2207 -17 2241 17
rect 2275 -17 2309 17
rect 2343 -17 2377 17
rect 2411 -17 2445 17
rect 2479 -17 2513 17
rect 2547 -17 2581 17
rect 2615 -17 2649 17
rect 2683 -17 2717 17
rect 2751 -17 2785 17
rect 2819 -17 2853 17
rect 2887 -17 2921 17
rect 2955 -17 2989 17
rect 3023 -17 3057 17
rect 3091 -17 3125 17
rect 3159 -17 3193 17
rect 3227 -17 3340 17
rect -1340 -40 3340 -17
rect -1340 -2240 -1300 -40
rect 3300 -2240 3340 -40
rect -1340 -2280 3340 -2240
<< nsubdiffcont >>
rect -1227 -17 -1193 17
rect -1159 -17 -1125 17
rect -1091 -17 -1057 17
rect -1023 -17 -989 17
rect -955 -17 -921 17
rect -887 -17 -853 17
rect -819 -17 -785 17
rect -751 -17 -717 17
rect -683 -17 -649 17
rect -615 -17 -581 17
rect -547 -17 -513 17
rect -479 -17 -445 17
rect -411 -17 -377 17
rect -343 -17 -309 17
rect -275 -17 -241 17
rect -207 -17 -173 17
rect -139 -17 -105 17
rect -71 -17 -37 17
rect -3 -17 31 17
rect 65 -17 99 17
rect 133 -17 167 17
rect 201 -17 235 17
rect 269 -17 303 17
rect 337 -17 371 17
rect 405 -17 439 17
rect 473 -17 507 17
rect 541 -17 575 17
rect 609 -17 643 17
rect 677 -17 711 17
rect 745 -17 779 17
rect 813 -17 847 17
rect 881 -17 915 17
rect 949 -17 983 17
rect 1017 -17 1051 17
rect 1085 -17 1119 17
rect 1153 -17 1187 17
rect 1221 -17 1255 17
rect 1289 -17 1323 17
rect 1357 -17 1391 17
rect 1425 -17 1459 17
rect 1493 -17 1527 17
rect 1561 -17 1595 17
rect 1629 -17 1663 17
rect 1697 -17 1731 17
rect 1765 -17 1799 17
rect 1833 -17 1867 17
rect 1901 -17 1935 17
rect 1969 -17 2003 17
rect 2037 -17 2071 17
rect 2105 -17 2139 17
rect 2173 -17 2207 17
rect 2241 -17 2275 17
rect 2309 -17 2343 17
rect 2377 -17 2411 17
rect 2445 -17 2479 17
rect 2513 -17 2547 17
rect 2581 -17 2615 17
rect 2649 -17 2683 17
rect 2717 -17 2751 17
rect 2785 -17 2819 17
rect 2853 -17 2887 17
rect 2921 -17 2955 17
rect 2989 -17 3023 17
rect 3057 -17 3091 17
rect 3125 -17 3159 17
rect 3193 -17 3227 17
<< locali >>
rect -1340 17 3340 40
rect -1340 -17 -1249 17
rect -1193 -17 -1177 17
rect -1125 -17 -1105 17
rect -1057 -17 -1033 17
rect -989 -17 -961 17
rect -921 -17 -889 17
rect -853 -17 -819 17
rect -783 -17 -751 17
rect -711 -17 -683 17
rect -639 -17 -615 17
rect -567 -17 -547 17
rect -495 -17 -479 17
rect -423 -17 -411 17
rect -351 -17 -343 17
rect -279 -17 -275 17
rect -173 -17 -169 17
rect -105 -17 -97 17
rect -37 -17 -25 17
rect 31 -17 47 17
rect 99 -17 119 17
rect 167 -17 191 17
rect 235 -17 263 17
rect 303 -17 335 17
rect 371 -17 405 17
rect 441 -17 473 17
rect 513 -17 541 17
rect 585 -17 609 17
rect 657 -17 677 17
rect 729 -17 745 17
rect 801 -17 813 17
rect 873 -17 881 17
rect 945 -17 949 17
rect 1051 -17 1055 17
rect 1119 -17 1127 17
rect 1187 -17 1199 17
rect 1255 -17 1271 17
rect 1323 -17 1343 17
rect 1391 -17 1415 17
rect 1459 -17 1487 17
rect 1527 -17 1559 17
rect 1595 -17 1629 17
rect 1665 -17 1697 17
rect 1737 -17 1765 17
rect 1809 -17 1833 17
rect 1881 -17 1901 17
rect 1953 -17 1969 17
rect 2025 -17 2037 17
rect 2097 -17 2105 17
rect 2169 -17 2173 17
rect 2275 -17 2279 17
rect 2343 -17 2351 17
rect 2411 -17 2423 17
rect 2479 -17 2495 17
rect 2547 -17 2567 17
rect 2615 -17 2639 17
rect 2683 -17 2711 17
rect 2751 -17 2783 17
rect 2819 -17 2853 17
rect 2889 -17 2921 17
rect 2961 -17 2989 17
rect 3033 -17 3057 17
rect 3105 -17 3125 17
rect 3177 -17 3193 17
rect 3249 -17 3340 17
rect -1340 -40 3340 -17
rect -1340 -2240 -1300 -40
rect 3300 -2240 3340 -40
rect -1340 -2280 3340 -2240
<< viali >>
rect -1249 -17 -1227 17
rect -1227 -17 -1215 17
rect -1177 -17 -1159 17
rect -1159 -17 -1143 17
rect -1105 -17 -1091 17
rect -1091 -17 -1071 17
rect -1033 -17 -1023 17
rect -1023 -17 -999 17
rect -961 -17 -955 17
rect -955 -17 -927 17
rect -889 -17 -887 17
rect -887 -17 -855 17
rect -817 -17 -785 17
rect -785 -17 -783 17
rect -745 -17 -717 17
rect -717 -17 -711 17
rect -673 -17 -649 17
rect -649 -17 -639 17
rect -601 -17 -581 17
rect -581 -17 -567 17
rect -529 -17 -513 17
rect -513 -17 -495 17
rect -457 -17 -445 17
rect -445 -17 -423 17
rect -385 -17 -377 17
rect -377 -17 -351 17
rect -313 -17 -309 17
rect -309 -17 -279 17
rect -241 -17 -207 17
rect -169 -17 -139 17
rect -139 -17 -135 17
rect -97 -17 -71 17
rect -71 -17 -63 17
rect -25 -17 -3 17
rect -3 -17 9 17
rect 47 -17 65 17
rect 65 -17 81 17
rect 119 -17 133 17
rect 133 -17 153 17
rect 191 -17 201 17
rect 201 -17 225 17
rect 263 -17 269 17
rect 269 -17 297 17
rect 335 -17 337 17
rect 337 -17 369 17
rect 407 -17 439 17
rect 439 -17 441 17
rect 479 -17 507 17
rect 507 -17 513 17
rect 551 -17 575 17
rect 575 -17 585 17
rect 623 -17 643 17
rect 643 -17 657 17
rect 695 -17 711 17
rect 711 -17 729 17
rect 767 -17 779 17
rect 779 -17 801 17
rect 839 -17 847 17
rect 847 -17 873 17
rect 911 -17 915 17
rect 915 -17 945 17
rect 983 -17 1017 17
rect 1055 -17 1085 17
rect 1085 -17 1089 17
rect 1127 -17 1153 17
rect 1153 -17 1161 17
rect 1199 -17 1221 17
rect 1221 -17 1233 17
rect 1271 -17 1289 17
rect 1289 -17 1305 17
rect 1343 -17 1357 17
rect 1357 -17 1377 17
rect 1415 -17 1425 17
rect 1425 -17 1449 17
rect 1487 -17 1493 17
rect 1493 -17 1521 17
rect 1559 -17 1561 17
rect 1561 -17 1593 17
rect 1631 -17 1663 17
rect 1663 -17 1665 17
rect 1703 -17 1731 17
rect 1731 -17 1737 17
rect 1775 -17 1799 17
rect 1799 -17 1809 17
rect 1847 -17 1867 17
rect 1867 -17 1881 17
rect 1919 -17 1935 17
rect 1935 -17 1953 17
rect 1991 -17 2003 17
rect 2003 -17 2025 17
rect 2063 -17 2071 17
rect 2071 -17 2097 17
rect 2135 -17 2139 17
rect 2139 -17 2169 17
rect 2207 -17 2241 17
rect 2279 -17 2309 17
rect 2309 -17 2313 17
rect 2351 -17 2377 17
rect 2377 -17 2385 17
rect 2423 -17 2445 17
rect 2445 -17 2457 17
rect 2495 -17 2513 17
rect 2513 -17 2529 17
rect 2567 -17 2581 17
rect 2581 -17 2601 17
rect 2639 -17 2649 17
rect 2649 -17 2673 17
rect 2711 -17 2717 17
rect 2717 -17 2745 17
rect 2783 -17 2785 17
rect 2785 -17 2817 17
rect 2855 -17 2887 17
rect 2887 -17 2889 17
rect 2927 -17 2955 17
rect 2955 -17 2961 17
rect 2999 -17 3023 17
rect 3023 -17 3033 17
rect 3071 -17 3091 17
rect 3091 -17 3105 17
rect 3143 -17 3159 17
rect 3159 -17 3177 17
rect 3215 -17 3227 17
rect 3227 -17 3249 17
<< metal1 >>
rect -1800 17 3340 40
rect -1800 -17 -1249 17
rect -1215 -17 -1177 17
rect -1143 -17 -1105 17
rect -1071 -17 -1033 17
rect -999 -17 -961 17
rect -927 -17 -889 17
rect -855 -17 -817 17
rect -783 -17 -745 17
rect -711 -17 -673 17
rect -639 -17 -601 17
rect -567 -17 -529 17
rect -495 -17 -457 17
rect -423 -17 -385 17
rect -351 -17 -313 17
rect -279 -17 -241 17
rect -207 -17 -169 17
rect -135 -17 -97 17
rect -63 -17 -25 17
rect 9 -17 47 17
rect 81 -17 119 17
rect 153 -17 191 17
rect 225 -17 263 17
rect 297 -17 335 17
rect 369 -17 407 17
rect 441 -17 479 17
rect 513 -17 551 17
rect 585 -17 623 17
rect 657 -17 695 17
rect 729 -17 767 17
rect 801 -17 839 17
rect 873 -17 911 17
rect 945 -17 983 17
rect 1017 -17 1055 17
rect 1089 -17 1127 17
rect 1161 -17 1199 17
rect 1233 -17 1271 17
rect 1305 -17 1343 17
rect 1377 -17 1415 17
rect 1449 -17 1487 17
rect 1521 -17 1559 17
rect 1593 -17 1631 17
rect 1665 -17 1703 17
rect 1737 -17 1775 17
rect 1809 -17 1847 17
rect 1881 -17 1919 17
rect 1953 -17 1991 17
rect 2025 -17 2063 17
rect 2097 -17 2135 17
rect 2169 -17 2207 17
rect 2241 -17 2279 17
rect 2313 -17 2351 17
rect 2385 -17 2423 17
rect 2457 -17 2495 17
rect 2529 -17 2567 17
rect 2601 -17 2639 17
rect 2673 -17 2711 17
rect 2745 -17 2783 17
rect 2817 -17 2855 17
rect 2889 -17 2927 17
rect 2961 -17 2999 17
rect 3033 -17 3071 17
rect 3105 -17 3143 17
rect 3177 -17 3215 17
rect 3249 -17 3340 17
rect -1800 -40 3340 -17
rect -1460 -137 -1380 -40
rect -1460 -189 -1446 -137
rect -1394 -189 -1380 -137
rect -1087 -134 -1010 -133
rect 620 -134 697 -133
rect -1087 -140 -1075 -134
rect -1460 -564 -1380 -189
rect -1140 -186 -1075 -140
rect -1023 -140 -1010 -134
rect -580 -135 -503 -134
rect -1023 -186 -840 -140
rect -580 -160 -568 -135
rect -1140 -200 -840 -186
rect -740 -187 -568 -160
rect -516 -160 -503 -135
rect 16 -135 93 -134
rect 16 -160 28 -135
rect -516 -187 -240 -160
rect -740 -200 -240 -187
rect -140 -187 28 -160
rect 80 -160 93 -135
rect 620 -160 632 -134
rect 80 -187 360 -160
rect -140 -200 360 -187
rect 460 -186 632 -160
rect 684 -160 697 -134
rect 2420 -136 2497 -135
rect 1823 -137 1900 -136
rect 1225 -138 1302 -137
rect 1225 -160 1237 -138
rect 684 -186 960 -160
rect 460 -200 960 -186
rect 1060 -190 1237 -160
rect 1289 -160 1302 -138
rect 1823 -140 1835 -137
rect 1289 -190 1560 -160
rect 1060 -200 1560 -190
rect 1660 -189 1835 -140
rect 1887 -140 1900 -137
rect 2420 -140 2432 -136
rect 1887 -189 2160 -140
rect 1660 -200 2160 -189
rect 2260 -188 2432 -140
rect 2484 -140 2497 -136
rect 2930 -136 3007 -135
rect 2930 -140 2942 -136
rect 2484 -188 2740 -140
rect 2260 -200 2740 -188
rect 2880 -188 2942 -140
rect 2994 -140 3007 -136
rect 2994 -188 3160 -140
rect 2880 -200 3160 -188
rect -900 -400 -840 -200
rect -1140 -460 -840 -400
rect -300 -420 -240 -200
rect 280 -400 360 -200
rect -740 -460 -240 -420
rect -140 -460 360 -400
rect 900 -420 960 -200
rect 1500 -400 1560 -200
rect 2080 -400 2160 -200
rect 2660 -400 2740 -200
rect 3100 -400 3160 -200
rect 480 -460 1440 -420
rect 1500 -459 1620 -440
rect 1500 -511 1536 -459
rect 1588 -511 1620 -459
rect 1700 -460 2160 -400
rect 2260 -460 2740 -400
rect 2880 -460 3160 -400
rect 1500 -560 1620 -511
rect -1462 -565 -1380 -564
rect -1462 -617 -1450 -565
rect -1398 -617 -1380 -565
rect -1460 -987 -1380 -617
rect -1120 -566 -840 -560
rect 20 -563 97 -562
rect -1120 -618 -1085 -566
rect -1033 -618 -840 -566
rect -567 -565 -490 -564
rect -567 -617 -555 -565
rect -503 -617 -490 -565
rect 20 -615 32 -563
rect 84 -615 97 -563
rect 1228 -564 1305 -563
rect 633 -565 710 -564
rect 633 -617 645 -565
rect 697 -617 710 -565
rect 1228 -616 1240 -564
rect 1292 -616 1305 -564
rect -1120 -620 -840 -618
rect -900 -820 -840 -620
rect -298 -693 -212 -678
rect -298 -745 -281 -693
rect -229 -745 -212 -693
rect -298 -759 -212 -745
rect 301 -698 387 -683
rect 301 -750 318 -698
rect 370 -750 387 -698
rect 301 -764 387 -750
rect 905 -701 991 -686
rect 905 -753 922 -701
rect 974 -753 991 -701
rect 905 -767 991 -753
rect 1500 -820 1580 -560
rect 2431 -561 2508 -560
rect 1824 -562 1901 -561
rect 1824 -614 1836 -562
rect 1888 -614 1901 -562
rect 2431 -613 2443 -561
rect 2495 -613 2508 -561
rect 2860 -561 3160 -560
rect 2860 -613 2937 -561
rect 2989 -613 3160 -561
rect 2860 -620 3160 -613
rect 2098 -696 2184 -681
rect 2098 -748 2115 -696
rect 2167 -748 2184 -696
rect 2098 -762 2184 -748
rect 2699 -696 2785 -681
rect 2699 -748 2716 -696
rect 2768 -748 2785 -696
rect 2699 -762 2785 -748
rect 3100 -820 3160 -620
rect -1140 -880 -840 -820
rect 441 -840 481 -835
rect -579 -843 -502 -842
rect -579 -895 -567 -843
rect -515 -895 -502 -843
rect 37 -846 114 -845
rect 37 -898 49 -846
rect 101 -898 114 -846
rect 380 -848 481 -840
rect 1815 -844 1892 -843
rect 379 -853 481 -848
rect 379 -905 394 -853
rect 446 -905 481 -853
rect 631 -849 708 -848
rect 631 -901 643 -849
rect 695 -901 708 -849
rect 1224 -849 1301 -848
rect 1224 -901 1236 -849
rect 1288 -901 1301 -849
rect 1815 -896 1827 -844
rect 1879 -896 1892 -844
rect 2422 -844 2499 -843
rect 2422 -896 2434 -844
rect 2486 -896 2499 -844
rect 2860 -880 3160 -820
rect 379 -910 481 -905
rect 380 -919 481 -910
rect 380 -920 458 -919
rect -1462 -988 -1380 -987
rect -1462 -1040 -1450 -988
rect -1398 -1040 -1380 -988
rect -1140 -986 -840 -980
rect -1140 -1038 -1059 -986
rect -1007 -1038 -840 -986
rect -568 -981 -491 -980
rect -568 -1033 -556 -981
rect -504 -1033 -491 -981
rect 26 -983 103 -982
rect 26 -1035 38 -983
rect 90 -1035 103 -983
rect -1140 -1040 -840 -1038
rect -1460 -1405 -1380 -1040
rect -900 -1240 -840 -1040
rect -303 -1121 -217 -1106
rect -303 -1173 -286 -1121
rect -234 -1173 -217 -1121
rect -303 -1187 -217 -1173
rect 272 -1114 350 -1102
rect 272 -1166 285 -1114
rect 337 -1166 350 -1114
rect 272 -1178 350 -1166
rect -1120 -1300 -840 -1240
rect -595 -1261 -518 -1260
rect -595 -1313 -583 -1261
rect -531 -1313 -518 -1261
rect 9 -1263 86 -1262
rect 9 -1315 21 -1263
rect 73 -1315 86 -1263
rect 380 -1279 420 -920
rect 637 -980 714 -979
rect 637 -1032 649 -980
rect 701 -1032 714 -980
rect 1235 -980 1312 -979
rect 1235 -1032 1247 -980
rect 1299 -1032 1312 -980
rect 1832 -980 1909 -979
rect 1832 -1032 1844 -980
rect 1896 -1032 1909 -980
rect 2434 -981 2511 -980
rect 2434 -1033 2446 -981
rect 2498 -1033 2511 -981
rect 2860 -981 3160 -980
rect 2860 -1033 2941 -981
rect 2993 -1033 3160 -981
rect 2860 -1040 3160 -1033
rect 895 -1116 981 -1101
rect 895 -1168 912 -1116
rect 964 -1168 981 -1116
rect 895 -1182 981 -1168
rect 1520 -1114 1620 -1040
rect 1520 -1166 1547 -1114
rect 1599 -1166 1620 -1114
rect 1520 -1240 1620 -1166
rect 2100 -1114 2186 -1099
rect 2100 -1166 2117 -1114
rect 2169 -1166 2186 -1114
rect 2100 -1180 2186 -1166
rect 2700 -1113 2786 -1098
rect 2700 -1165 2717 -1113
rect 2769 -1165 2786 -1113
rect 2700 -1179 2786 -1165
rect 3100 -1240 3160 -1040
rect 627 -1265 704 -1264
rect 353 -1280 430 -1279
rect 353 -1332 365 -1280
rect 417 -1332 430 -1280
rect 627 -1317 639 -1265
rect 691 -1317 704 -1265
rect 1062 -1286 1460 -1246
rect 362 -1337 422 -1332
rect -1460 -1457 -1445 -1405
rect -1393 -1457 -1380 -1405
rect -1460 -2117 -1380 -1457
rect -1140 -1402 -860 -1400
rect -1140 -1454 -1070 -1402
rect -1018 -1454 -860 -1402
rect -1140 -1460 -860 -1454
rect -572 -1403 -495 -1402
rect -572 -1455 -560 -1403
rect -508 -1455 -495 -1403
rect 27 -1403 104 -1402
rect 27 -1455 39 -1403
rect 91 -1455 104 -1403
rect -920 -1660 -860 -1460
rect -299 -1540 -213 -1525
rect -299 -1592 -282 -1540
rect -230 -1592 -213 -1540
rect 272 -1535 349 -1534
rect 272 -1587 284 -1535
rect 336 -1587 349 -1535
rect -299 -1606 -213 -1592
rect -1140 -1720 -860 -1660
rect 380 -1680 420 -1337
rect 1062 -1338 1196 -1286
rect 1248 -1338 1260 -1286
rect 1312 -1338 1460 -1286
rect 1825 -1259 1902 -1258
rect 1825 -1311 1837 -1259
rect 1889 -1311 1902 -1259
rect 2432 -1263 2509 -1262
rect 2432 -1315 2444 -1263
rect 2496 -1315 2509 -1263
rect 2860 -1300 3160 -1240
rect 3220 -1267 3300 -560
rect 3380 -849 3460 -560
rect 3380 -901 3395 -849
rect 3447 -901 3460 -849
rect 3380 -1258 3460 -901
rect 3220 -1268 3307 -1267
rect 1062 -1340 1460 -1338
rect 3220 -1320 3242 -1268
rect 3294 -1320 3307 -1268
rect 1180 -1349 1328 -1340
rect 626 -1400 703 -1399
rect 626 -1452 638 -1400
rect 690 -1452 703 -1400
rect 1231 -1402 1308 -1401
rect 1231 -1454 1243 -1402
rect 1295 -1454 1308 -1402
rect 2428 -1402 2505 -1401
rect 1827 -1404 1904 -1403
rect 1827 -1456 1839 -1404
rect 1891 -1456 1904 -1404
rect 2428 -1454 2440 -1402
rect 2492 -1454 2505 -1402
rect 2860 -1402 3160 -1400
rect 2860 -1454 2944 -1402
rect 2996 -1454 3160 -1402
rect 2860 -1460 3160 -1454
rect 907 -1539 993 -1524
rect 907 -1591 924 -1539
rect 976 -1591 993 -1539
rect 907 -1605 993 -1591
rect 1504 -1539 1590 -1524
rect 1504 -1591 1521 -1539
rect 1573 -1591 1590 -1539
rect 1504 -1605 1590 -1591
rect 2094 -1544 2180 -1529
rect 2094 -1596 2111 -1544
rect 2163 -1596 2180 -1544
rect 2094 -1610 2180 -1596
rect 2704 -1539 2790 -1524
rect 2704 -1591 2721 -1539
rect 2773 -1591 2790 -1539
rect 2704 -1605 2790 -1591
rect 3100 -1660 3160 -1460
rect 31 -1683 108 -1682
rect -581 -1684 -504 -1683
rect -581 -1736 -569 -1684
rect -517 -1736 -504 -1684
rect 31 -1735 43 -1683
rect 95 -1735 108 -1683
rect 380 -1684 479 -1680
rect 1823 -1684 1900 -1683
rect 380 -1690 502 -1684
rect 379 -1695 502 -1690
rect 379 -1747 394 -1695
rect 446 -1747 502 -1695
rect 597 -1690 674 -1689
rect 597 -1742 609 -1690
rect 661 -1742 674 -1690
rect 1214 -1690 1291 -1689
rect 1214 -1742 1226 -1690
rect 1278 -1742 1291 -1690
rect 1823 -1736 1835 -1684
rect 1887 -1736 1900 -1684
rect 2429 -1684 2506 -1683
rect 2429 -1736 2441 -1684
rect 2493 -1736 2506 -1684
rect 2880 -1720 3160 -1660
rect 379 -1752 502 -1747
rect 380 -1760 502 -1752
rect -1140 -1880 -860 -1840
rect -740 -1880 -260 -1820
rect -140 -1880 320 -1820
rect -940 -2100 -860 -1880
rect -320 -2080 -260 -1880
rect 260 -2080 320 -1880
rect -1460 -2169 -1447 -2117
rect -1395 -2169 -1380 -2117
rect -1140 -2108 -860 -2100
rect -1140 -2140 -1078 -2108
rect -1090 -2160 -1078 -2140
rect -1026 -2140 -860 -2108
rect -740 -2108 -260 -2080
rect -740 -2140 -558 -2108
rect -1026 -2160 -1013 -2140
rect -570 -2160 -558 -2140
rect -506 -2140 -260 -2108
rect -140 -2108 320 -2080
rect -140 -2140 22 -2108
rect -506 -2160 -493 -2140
rect 10 -2160 22 -2140
rect 74 -2140 320 -2108
rect 74 -2160 87 -2140
rect -1460 -2180 -1380 -2169
rect 380 -2320 420 -1760
rect 458 -1761 502 -1760
rect 2860 -1840 3120 -1820
rect 460 -1880 940 -1840
rect 1060 -1880 1540 -1840
rect 1660 -1880 2140 -1840
rect 2260 -1880 2740 -1840
rect 2860 -1880 3140 -1840
rect 860 -2080 940 -1880
rect 1480 -2080 1540 -1880
rect 2060 -2080 2140 -1880
rect 2680 -2080 2740 -1880
rect 3080 -2080 3140 -1880
rect 480 -2108 940 -2080
rect 480 -2140 622 -2108
rect 610 -2160 622 -2140
rect 674 -2140 940 -2108
rect 1060 -2108 1540 -2080
rect 1060 -2140 1242 -2108
rect 674 -2160 687 -2140
rect 1230 -2160 1242 -2140
rect 1294 -2140 1540 -2108
rect 1660 -2108 2140 -2080
rect 1660 -2140 1822 -2108
rect 1294 -2160 1307 -2140
rect 1810 -2160 1822 -2140
rect 1874 -2140 2140 -2108
rect 2260 -2108 2740 -2080
rect 2260 -2140 2422 -2108
rect 1874 -2160 1887 -2140
rect 2410 -2160 2422 -2140
rect 2474 -2140 2740 -2108
rect 2860 -2108 3140 -2080
rect 2860 -2140 2942 -2108
rect 2474 -2160 2487 -2140
rect 2912 -2150 2942 -2140
rect 2930 -2160 2942 -2150
rect 2994 -2140 3140 -2108
rect 2994 -2160 3007 -2140
rect 380 -2337 460 -2320
rect 380 -2389 392 -2337
rect 444 -2389 460 -2337
rect 380 -2400 460 -2389
rect 3220 -2340 3300 -1320
rect 3220 -2392 3236 -2340
rect 3288 -2392 3300 -2340
rect 3220 -2400 3300 -2392
rect 3380 -1335 3461 -1258
rect 3380 -1387 3392 -1335
rect 3444 -1387 3461 -1335
rect 3380 -1401 3461 -1387
rect 3380 -1676 3460 -1401
rect 3380 -1728 3393 -1676
rect 3445 -1728 3460 -1676
rect 3380 -2446 3460 -1728
rect 3380 -2498 3395 -2446
rect 3447 -2498 3460 -2446
rect 3380 -2510 3460 -2498
<< via1 >>
rect -1446 -189 -1394 -137
rect -1075 -186 -1023 -134
rect -568 -187 -516 -135
rect 28 -187 80 -135
rect 632 -186 684 -134
rect 1237 -190 1289 -138
rect 1835 -189 1887 -137
rect 2432 -188 2484 -136
rect 2942 -188 2994 -136
rect 1536 -511 1588 -459
rect -1450 -617 -1398 -565
rect -1085 -618 -1033 -566
rect -555 -617 -503 -565
rect 32 -615 84 -563
rect 645 -617 697 -565
rect 1240 -616 1292 -564
rect -281 -745 -229 -693
rect 318 -750 370 -698
rect 922 -753 974 -701
rect 1836 -614 1888 -562
rect 2443 -613 2495 -561
rect 2937 -613 2989 -561
rect 2115 -748 2167 -696
rect 2716 -748 2768 -696
rect -567 -895 -515 -843
rect 49 -898 101 -846
rect 394 -905 446 -853
rect 643 -901 695 -849
rect 1236 -901 1288 -849
rect 1827 -896 1879 -844
rect 2434 -896 2486 -844
rect -1450 -1040 -1398 -988
rect -1059 -1038 -1007 -986
rect -556 -1033 -504 -981
rect 38 -1035 90 -983
rect -286 -1173 -234 -1121
rect 285 -1166 337 -1114
rect -583 -1313 -531 -1261
rect 21 -1315 73 -1263
rect 649 -1032 701 -980
rect 1247 -1032 1299 -980
rect 1844 -1032 1896 -980
rect 2446 -1033 2498 -981
rect 2941 -1033 2993 -981
rect 912 -1168 964 -1116
rect 1547 -1166 1599 -1114
rect 2117 -1166 2169 -1114
rect 2717 -1165 2769 -1113
rect 365 -1332 417 -1280
rect 639 -1317 691 -1265
rect -1445 -1457 -1393 -1405
rect -1070 -1454 -1018 -1402
rect -560 -1455 -508 -1403
rect 39 -1455 91 -1403
rect -282 -1592 -230 -1540
rect 284 -1587 336 -1535
rect 1196 -1338 1248 -1286
rect 1260 -1338 1312 -1286
rect 1837 -1311 1889 -1259
rect 2444 -1315 2496 -1263
rect 3395 -901 3447 -849
rect 3242 -1320 3294 -1268
rect 638 -1452 690 -1400
rect 1243 -1454 1295 -1402
rect 1839 -1456 1891 -1404
rect 2440 -1454 2492 -1402
rect 2944 -1454 2996 -1402
rect 924 -1591 976 -1539
rect 1521 -1591 1573 -1539
rect 2111 -1596 2163 -1544
rect 2721 -1591 2773 -1539
rect -569 -1736 -517 -1684
rect 43 -1735 95 -1683
rect 394 -1747 446 -1695
rect 609 -1742 661 -1690
rect 1226 -1742 1278 -1690
rect 1835 -1736 1887 -1684
rect 2441 -1736 2493 -1684
rect -1447 -2169 -1395 -2117
rect -1078 -2160 -1026 -2108
rect -558 -2160 -506 -2108
rect 22 -2160 74 -2108
rect 622 -2160 674 -2108
rect 1242 -2160 1294 -2108
rect 1822 -2160 1874 -2108
rect 2422 -2160 2474 -2108
rect 2942 -2160 2994 -2108
rect 392 -2389 444 -2337
rect 3236 -2392 3288 -2340
rect 3392 -1387 3444 -1335
rect 3393 -1728 3445 -1676
rect 3395 -2498 3447 -2446
<< metal2 >>
rect -1460 -134 3060 -120
rect -1460 -137 -1075 -134
rect -1460 -189 -1446 -137
rect -1394 -186 -1075 -137
rect -1023 -135 632 -134
rect -1023 -186 -568 -135
rect -1394 -187 -568 -186
rect -516 -187 28 -135
rect 80 -186 632 -135
rect 684 -136 3060 -134
rect 684 -137 2432 -136
rect 684 -138 1835 -137
rect 684 -186 1237 -138
rect 80 -187 1237 -186
rect -1394 -189 1237 -187
rect -1460 -190 1237 -189
rect 1289 -189 1835 -138
rect 1887 -188 2432 -137
rect 2484 -188 2942 -136
rect 2994 -188 3060 -136
rect 1887 -189 3060 -188
rect 1289 -190 3060 -189
rect -1460 -200 3060 -190
rect 1518 -457 1607 -439
rect 1518 -513 1534 -457
rect 1590 -513 1607 -457
rect 1518 -531 1607 -513
rect -1461 -560 -1380 -540
rect -557 -560 -500 -554
rect 30 -560 87 -552
rect 643 -560 700 -554
rect 1238 -560 1295 -553
rect 1834 -560 1891 -551
rect 2441 -560 2498 -550
rect 2935 -560 2992 -550
rect -1461 -561 3080 -560
rect -1461 -562 2443 -561
rect -1461 -563 1836 -562
rect -1461 -565 32 -563
rect -1461 -617 -1450 -565
rect -1398 -566 -555 -565
rect -1398 -617 -1085 -566
rect -1461 -618 -1085 -617
rect -1033 -617 -555 -566
rect -503 -615 32 -565
rect 84 -564 1836 -563
rect 84 -565 1240 -564
rect 84 -615 645 -565
rect -503 -617 645 -615
rect 697 -616 1240 -565
rect 1292 -614 1836 -564
rect 1888 -613 2443 -562
rect 2495 -613 2937 -561
rect 2989 -613 3080 -561
rect 1888 -614 3080 -613
rect 1292 -616 3080 -614
rect 697 -617 3080 -616
rect -1033 -618 3080 -617
rect -1461 -620 3080 -618
rect -1461 -641 -1380 -620
rect -557 -627 -500 -620
rect 30 -625 87 -620
rect 643 -627 700 -620
rect 1238 -626 1295 -620
rect 1834 -624 1891 -620
rect 2441 -623 2498 -620
rect 2935 -623 2992 -620
rect -288 -691 -222 -668
rect -288 -747 -283 -691
rect -227 -747 -222 -691
rect -288 -769 -222 -747
rect 311 -696 377 -673
rect 311 -752 316 -696
rect 372 -752 377 -696
rect 311 -774 377 -752
rect 915 -699 981 -676
rect 915 -755 920 -699
rect 976 -755 981 -699
rect 915 -777 981 -755
rect 2108 -694 2174 -671
rect 2108 -750 2113 -694
rect 2169 -750 2174 -694
rect 2108 -772 2174 -750
rect 2709 -694 2775 -671
rect 2709 -750 2714 -694
rect 2770 -750 2775 -694
rect 2709 -772 2775 -750
rect -820 -840 -760 -828
rect -569 -840 -512 -832
rect 47 -840 104 -835
rect 389 -840 452 -838
rect 641 -840 698 -838
rect 1234 -840 1291 -838
rect 1680 -840 1760 -838
rect 1825 -840 1882 -833
rect 2432 -840 2489 -833
rect 3393 -840 3450 -838
rect -820 -841 260 -840
rect -820 -897 -818 -841
rect -762 -843 260 -841
rect -762 -895 -567 -843
rect -515 -846 260 -843
rect -515 -895 49 -846
rect -762 -897 49 -895
rect -820 -898 49 -897
rect 101 -898 260 -846
rect -820 -900 260 -898
rect 380 -849 1460 -840
rect 380 -853 643 -849
rect -820 -910 -760 -900
rect -569 -905 -512 -900
rect 47 -908 104 -900
rect 380 -905 394 -853
rect 446 -901 643 -853
rect 695 -901 1236 -849
rect 1288 -901 1460 -849
rect 1680 -844 3460 -840
rect 1680 -896 1827 -844
rect 1879 -896 2434 -844
rect 2486 -849 3460 -844
rect 2486 -896 3395 -849
rect 1680 -900 3395 -896
rect 446 -905 1460 -901
rect 380 -920 1460 -905
rect 1825 -906 1882 -900
rect 2432 -906 2489 -900
rect 3393 -901 3395 -900
rect 3447 -900 3460 -849
rect 3447 -901 3450 -900
rect 3393 -911 3450 -901
rect -1460 -980 -1379 -959
rect -1061 -980 -1004 -975
rect -558 -980 -501 -970
rect 36 -980 93 -972
rect 647 -980 704 -969
rect 1245 -980 1302 -969
rect 1842 -980 1899 -969
rect 2444 -980 2501 -970
rect 2939 -980 2996 -970
rect -1460 -981 649 -980
rect -1460 -986 -556 -981
rect -1460 -988 -1059 -986
rect -1460 -1040 -1450 -988
rect -1398 -1038 -1059 -988
rect -1007 -1033 -556 -986
rect -504 -983 649 -981
rect -504 -1033 38 -983
rect -1007 -1035 38 -1033
rect 90 -1032 649 -983
rect 701 -1032 1247 -980
rect 1299 -1032 1844 -980
rect 1896 -981 3080 -980
rect 1896 -1032 2446 -981
rect 90 -1033 2446 -1032
rect 2498 -1033 2941 -981
rect 2993 -1033 3080 -981
rect 90 -1035 3080 -1033
rect -1007 -1038 3080 -1035
rect -1398 -1040 3080 -1038
rect -1460 -1060 -1379 -1040
rect -1061 -1048 -1004 -1040
rect -558 -1043 -501 -1040
rect 36 -1045 93 -1040
rect 647 -1042 704 -1040
rect 1245 -1042 1302 -1040
rect 1842 -1042 1899 -1040
rect 2444 -1043 2501 -1040
rect 2939 -1043 2996 -1040
rect -293 -1119 -227 -1096
rect -293 -1175 -288 -1119
rect -232 -1175 -227 -1119
rect -293 -1197 -227 -1175
rect 282 -1112 340 -1092
rect 282 -1168 283 -1112
rect 339 -1168 340 -1112
rect 282 -1188 340 -1168
rect 905 -1114 971 -1091
rect 905 -1170 910 -1114
rect 966 -1170 971 -1114
rect 905 -1192 971 -1170
rect 1540 -1112 1606 -1089
rect 1540 -1168 1545 -1112
rect 1601 -1168 1606 -1112
rect 1540 -1190 1606 -1168
rect 2110 -1112 2176 -1089
rect 2110 -1168 2115 -1112
rect 2171 -1168 2176 -1112
rect 2110 -1190 2176 -1168
rect 2710 -1111 2776 -1088
rect 2710 -1167 2715 -1111
rect 2771 -1167 2776 -1111
rect 2710 -1189 2776 -1167
rect -585 -1260 -528 -1250
rect 19 -1260 76 -1252
rect 637 -1260 694 -1254
rect 1835 -1259 1892 -1248
rect 1835 -1260 1837 -1259
rect -740 -1261 860 -1260
rect -740 -1313 -583 -1261
rect -531 -1263 860 -1261
rect -531 -1313 21 -1263
rect -740 -1315 21 -1313
rect 73 -1265 860 -1263
rect 73 -1280 639 -1265
rect 73 -1315 365 -1280
rect -740 -1320 365 -1315
rect -585 -1323 -528 -1320
rect 19 -1325 76 -1320
rect 339 -1332 365 -1320
rect 417 -1317 639 -1280
rect 691 -1317 860 -1265
rect 417 -1320 860 -1317
rect 1190 -1284 1318 -1265
rect 1190 -1286 1226 -1284
rect 1282 -1286 1318 -1284
rect 417 -1332 421 -1320
rect 637 -1327 694 -1320
rect 339 -1341 421 -1332
rect 1190 -1338 1196 -1286
rect 1312 -1338 1318 -1286
rect 1800 -1311 1837 -1260
rect 1889 -1260 1892 -1259
rect 2442 -1260 2499 -1252
rect 3240 -1260 3297 -1257
rect 1889 -1263 3300 -1260
rect 1889 -1311 2444 -1263
rect 1800 -1315 2444 -1311
rect 2496 -1268 3300 -1263
rect 2496 -1315 3242 -1268
rect 1800 -1320 3242 -1315
rect 3294 -1320 3300 -1268
rect 1835 -1321 1892 -1320
rect 2442 -1325 2499 -1320
rect 3240 -1330 3297 -1320
rect 1190 -1340 1226 -1338
rect 1282 -1340 1318 -1338
rect 363 -1342 420 -1341
rect 1190 -1359 1318 -1340
rect 3385 -1333 3451 -1310
rect -1460 -1400 -1379 -1379
rect 3385 -1389 3390 -1333
rect 3446 -1389 3451 -1333
rect -1072 -1400 -1015 -1391
rect -562 -1400 -505 -1392
rect 37 -1400 94 -1392
rect 636 -1400 693 -1389
rect 1241 -1400 1298 -1391
rect 1837 -1400 1894 -1393
rect 2438 -1400 2495 -1391
rect 2942 -1400 2999 -1391
rect -1460 -1402 638 -1400
rect -1460 -1405 -1070 -1402
rect -1460 -1457 -1445 -1405
rect -1393 -1454 -1070 -1405
rect -1018 -1403 638 -1402
rect -1018 -1454 -560 -1403
rect -1393 -1455 -560 -1454
rect -508 -1455 39 -1403
rect 91 -1452 638 -1403
rect 690 -1402 3080 -1400
rect 690 -1452 1243 -1402
rect 91 -1454 1243 -1452
rect 1295 -1404 2440 -1402
rect 1295 -1454 1839 -1404
rect 91 -1455 1839 -1454
rect -1393 -1456 1839 -1455
rect 1891 -1454 2440 -1404
rect 2492 -1454 2944 -1402
rect 2996 -1454 3080 -1402
rect 3385 -1411 3451 -1389
rect 1891 -1456 3080 -1454
rect -1393 -1457 3080 -1456
rect -1460 -1460 3080 -1457
rect -1460 -1480 -1379 -1460
rect -1072 -1464 -1015 -1460
rect -562 -1465 -505 -1460
rect 37 -1465 94 -1460
rect 636 -1462 693 -1460
rect 1241 -1464 1298 -1460
rect 1837 -1466 1894 -1460
rect 2438 -1464 2495 -1460
rect 2942 -1464 2999 -1460
rect -289 -1538 -223 -1515
rect 284 -1524 340 -1518
rect -289 -1594 -284 -1538
rect -228 -1594 -223 -1538
rect -289 -1616 -223 -1594
rect 282 -1534 340 -1524
rect 282 -1590 284 -1534
rect 282 -1597 340 -1590
rect 284 -1605 340 -1597
rect 917 -1537 983 -1514
rect 917 -1593 922 -1537
rect 978 -1593 983 -1537
rect 917 -1615 983 -1593
rect 1514 -1537 1580 -1514
rect 1514 -1593 1519 -1537
rect 1575 -1593 1580 -1537
rect 1514 -1615 1580 -1593
rect 2104 -1542 2170 -1519
rect 2104 -1598 2109 -1542
rect 2165 -1598 2170 -1542
rect 2104 -1620 2170 -1598
rect 2714 -1537 2780 -1514
rect 2714 -1593 2719 -1537
rect 2775 -1593 2780 -1537
rect 2714 -1615 2780 -1593
rect -820 -1680 -760 -1668
rect -571 -1680 -514 -1673
rect 41 -1680 98 -1672
rect 607 -1680 664 -1679
rect 1224 -1680 1281 -1679
rect 1600 -1680 1660 -1668
rect 1833 -1680 1890 -1673
rect 2439 -1680 2496 -1673
rect 3391 -1676 3448 -1665
rect 3391 -1680 3393 -1676
rect -820 -1681 260 -1680
rect -820 -1737 -818 -1681
rect -762 -1683 260 -1681
rect -762 -1684 43 -1683
rect -762 -1736 -569 -1684
rect -517 -1735 43 -1684
rect 95 -1735 260 -1683
rect -517 -1736 260 -1735
rect -762 -1737 260 -1736
rect -820 -1740 260 -1737
rect 380 -1690 1460 -1680
rect 380 -1695 609 -1690
rect -820 -1750 -760 -1740
rect -571 -1746 -514 -1740
rect 41 -1745 98 -1740
rect 380 -1747 394 -1695
rect 446 -1742 609 -1695
rect 661 -1742 1226 -1690
rect 1278 -1742 1460 -1690
rect 446 -1747 1460 -1742
rect 380 -1760 1460 -1747
rect 1600 -1684 3393 -1680
rect 1600 -1736 1835 -1684
rect 1887 -1736 2441 -1684
rect 2493 -1728 3393 -1684
rect 3445 -1680 3448 -1676
rect 3445 -1728 3460 -1680
rect 2493 -1736 3460 -1728
rect 1600 -1740 3460 -1736
rect 1600 -1750 1660 -1740
rect 1833 -1746 1890 -1740
rect 2439 -1746 2496 -1740
rect 389 -1762 452 -1760
rect -1080 -2100 -1023 -2097
rect -560 -2100 -503 -2097
rect 20 -2100 77 -2097
rect 620 -2100 677 -2097
rect 1240 -2100 1297 -2097
rect 1820 -2100 1877 -2097
rect 2420 -2100 2477 -2097
rect 2940 -2100 2997 -2097
rect -1460 -2108 3140 -2100
rect -1460 -2117 -1078 -2108
rect -1460 -2169 -1447 -2117
rect -1395 -2160 -1078 -2117
rect -1026 -2160 -558 -2108
rect -506 -2160 22 -2108
rect 74 -2160 622 -2108
rect 674 -2160 1242 -2108
rect 1294 -2160 1822 -2108
rect 1874 -2160 2422 -2108
rect 2474 -2160 2942 -2108
rect 2994 -2160 3140 -2108
rect -1395 -2169 3140 -2160
rect -1460 -2180 3140 -2169
rect 380 -2337 3300 -2320
rect 380 -2389 392 -2337
rect 444 -2340 3300 -2337
rect 444 -2389 3236 -2340
rect 380 -2392 3236 -2389
rect 3288 -2392 3300 -2340
rect 380 -2400 3300 -2392
rect 3234 -2402 3291 -2400
rect -820 -2443 3460 -2430
rect -820 -2499 -810 -2443
rect -754 -2446 3460 -2443
rect -754 -2498 3395 -2446
rect 3447 -2498 3460 -2446
rect -754 -2499 3460 -2498
rect -820 -2510 3460 -2499
<< via2 >>
rect 1534 -459 1590 -457
rect 1534 -511 1536 -459
rect 1536 -511 1588 -459
rect 1588 -511 1590 -459
rect 1534 -513 1590 -511
rect -283 -693 -227 -691
rect -283 -745 -281 -693
rect -281 -745 -229 -693
rect -229 -745 -227 -693
rect -283 -747 -227 -745
rect 316 -698 372 -696
rect 316 -750 318 -698
rect 318 -750 370 -698
rect 370 -750 372 -698
rect 316 -752 372 -750
rect 920 -701 976 -699
rect 920 -753 922 -701
rect 922 -753 974 -701
rect 974 -753 976 -701
rect 920 -755 976 -753
rect 2113 -696 2169 -694
rect 2113 -748 2115 -696
rect 2115 -748 2167 -696
rect 2167 -748 2169 -696
rect 2113 -750 2169 -748
rect 2714 -696 2770 -694
rect 2714 -748 2716 -696
rect 2716 -748 2768 -696
rect 2768 -748 2770 -696
rect 2714 -750 2770 -748
rect -818 -897 -762 -841
rect -288 -1121 -232 -1119
rect -288 -1173 -286 -1121
rect -286 -1173 -234 -1121
rect -234 -1173 -232 -1121
rect -288 -1175 -232 -1173
rect 283 -1114 339 -1112
rect 283 -1166 285 -1114
rect 285 -1166 337 -1114
rect 337 -1166 339 -1114
rect 283 -1168 339 -1166
rect 910 -1116 966 -1114
rect 910 -1168 912 -1116
rect 912 -1168 964 -1116
rect 964 -1168 966 -1116
rect 910 -1170 966 -1168
rect 1545 -1114 1601 -1112
rect 1545 -1166 1547 -1114
rect 1547 -1166 1599 -1114
rect 1599 -1166 1601 -1114
rect 1545 -1168 1601 -1166
rect 2115 -1114 2171 -1112
rect 2115 -1166 2117 -1114
rect 2117 -1166 2169 -1114
rect 2169 -1166 2171 -1114
rect 2115 -1168 2171 -1166
rect 2715 -1113 2771 -1111
rect 2715 -1165 2717 -1113
rect 2717 -1165 2769 -1113
rect 2769 -1165 2771 -1113
rect 2715 -1167 2771 -1165
rect 1226 -1286 1282 -1284
rect 1226 -1338 1248 -1286
rect 1248 -1338 1260 -1286
rect 1260 -1338 1282 -1286
rect 1226 -1340 1282 -1338
rect 3390 -1335 3446 -1333
rect 3390 -1387 3392 -1335
rect 3392 -1387 3444 -1335
rect 3444 -1387 3446 -1335
rect 3390 -1389 3446 -1387
rect -284 -1540 -228 -1538
rect -284 -1592 -282 -1540
rect -282 -1592 -230 -1540
rect -230 -1592 -228 -1540
rect -284 -1594 -228 -1592
rect 284 -1535 340 -1534
rect 284 -1587 336 -1535
rect 336 -1587 340 -1535
rect 284 -1590 340 -1587
rect 922 -1539 978 -1537
rect 922 -1591 924 -1539
rect 924 -1591 976 -1539
rect 976 -1591 978 -1539
rect 922 -1593 978 -1591
rect 1519 -1539 1575 -1537
rect 1519 -1591 1521 -1539
rect 1521 -1591 1573 -1539
rect 1573 -1591 1575 -1539
rect 1519 -1593 1575 -1591
rect 2109 -1544 2165 -1542
rect 2109 -1596 2111 -1544
rect 2111 -1596 2163 -1544
rect 2163 -1596 2165 -1544
rect 2109 -1598 2165 -1596
rect 2719 -1539 2775 -1537
rect 2719 -1591 2721 -1539
rect 2721 -1591 2773 -1539
rect 2773 -1591 2775 -1539
rect 2719 -1593 2775 -1591
rect -818 -1737 -762 -1681
rect -810 -2499 -754 -2443
<< metal3 >>
rect 1508 -453 1617 -444
rect 1508 -480 1530 -453
rect 900 -486 1019 -480
rect 900 -550 926 -486
rect 990 -550 1019 -486
rect 900 -560 1019 -550
rect 1500 -517 1530 -480
rect 1594 -517 1617 -453
rect 1500 -526 1617 -517
rect -300 -673 -220 -660
rect -300 -687 -212 -673
rect -300 -751 -287 -687
rect -223 -751 -212 -687
rect -300 -764 -212 -751
rect 300 -678 380 -660
rect 300 -692 387 -678
rect 300 -756 312 -692
rect 376 -756 387 -692
rect -300 -780 -220 -764
rect 300 -769 387 -756
rect 900 -681 980 -560
rect 1500 -600 1580 -526
rect 2100 -676 2180 -660
rect 2700 -676 2780 -660
rect 1550 -680 1636 -679
rect 900 -699 991 -681
rect 900 -755 920 -699
rect 976 -755 991 -699
rect 300 -780 380 -769
rect 900 -772 991 -755
rect 1540 -688 1636 -680
rect 1540 -752 1561 -688
rect 1625 -752 1636 -688
rect 1540 -760 1636 -752
rect 2098 -690 2184 -676
rect 2098 -754 2109 -690
rect 2173 -754 2184 -690
rect -830 -841 -750 -833
rect -830 -897 -818 -841
rect -762 -897 -750 -841
rect -830 -905 -750 -897
rect -820 -1673 -760 -905
rect -320 -1101 -240 -1080
rect 300 -1097 380 -1080
rect 900 -1096 980 -772
rect 1540 -1094 1620 -760
rect 2098 -767 2184 -754
rect 2699 -690 2785 -676
rect 2699 -754 2710 -690
rect 2774 -754 2785 -690
rect 2699 -767 2785 -754
rect 2100 -780 2180 -767
rect 2700 -780 2780 -767
rect -320 -1115 -217 -1101
rect -320 -1179 -292 -1115
rect -228 -1179 -217 -1115
rect 267 -1106 380 -1097
rect 267 -1170 278 -1106
rect 342 -1170 380 -1106
rect 267 -1178 380 -1170
rect -320 -1192 -217 -1179
rect 272 -1183 380 -1178
rect -320 -1200 -240 -1192
rect 300 -1200 380 -1183
rect 895 -1110 981 -1096
rect 895 -1174 906 -1110
rect 970 -1174 981 -1110
rect 895 -1187 981 -1174
rect 1530 -1112 1620 -1094
rect 1530 -1168 1545 -1112
rect 1601 -1168 1620 -1112
rect 1530 -1185 1620 -1168
rect -300 -1520 -220 -1500
rect 280 -1519 360 -1500
rect -300 -1534 -213 -1520
rect -300 -1598 -288 -1534
rect -224 -1598 -213 -1534
rect -300 -1611 -213 -1598
rect 270 -1528 360 -1519
rect 270 -1592 281 -1528
rect 345 -1592 360 -1528
rect 270 -1600 360 -1592
rect -300 -1620 -220 -1611
rect 280 -1620 360 -1600
rect 900 -1519 980 -1187
rect 1540 -1240 1620 -1185
rect 2080 -1094 2160 -1080
rect 2700 -1093 2780 -1080
rect 2080 -1108 2186 -1094
rect 2080 -1172 2111 -1108
rect 2175 -1172 2186 -1108
rect 2080 -1185 2186 -1172
rect 2700 -1107 2786 -1093
rect 2700 -1171 2711 -1107
rect 2775 -1171 2786 -1107
rect 2700 -1184 2786 -1171
rect 2080 -1200 2160 -1185
rect 2700 -1200 2780 -1184
rect 1180 -1280 1328 -1270
rect 1180 -1344 1222 -1280
rect 1286 -1344 1328 -1280
rect 3380 -1315 3460 -1300
rect 1180 -1354 1328 -1344
rect 3375 -1329 3461 -1315
rect 3375 -1393 3386 -1329
rect 3450 -1393 3461 -1329
rect 3375 -1406 3461 -1393
rect 3380 -1420 3460 -1406
rect 1500 -1519 1580 -1500
rect 900 -1537 993 -1519
rect 900 -1593 922 -1537
rect 978 -1593 993 -1537
rect 900 -1610 993 -1593
rect 1500 -1537 1590 -1519
rect 2100 -1524 2180 -1500
rect 1500 -1593 1519 -1537
rect 1575 -1593 1590 -1537
rect 1500 -1610 1590 -1593
rect 2094 -1538 2180 -1524
rect 2094 -1602 2105 -1538
rect 2169 -1602 2180 -1538
rect -830 -1681 -750 -1673
rect -830 -1737 -818 -1681
rect -762 -1737 -750 -1681
rect -830 -1745 -750 -1737
rect -820 -2430 -760 -1745
rect 900 -1751 980 -1610
rect 1500 -1745 1580 -1610
rect 2094 -1615 2180 -1602
rect 2100 -1620 2180 -1615
rect 2700 -1519 2780 -1500
rect 2700 -1533 2790 -1519
rect 2700 -1597 2715 -1533
rect 2779 -1597 2790 -1533
rect 2700 -1610 2790 -1597
rect 2700 -1620 2780 -1610
rect 1493 -1747 1584 -1745
rect 896 -1753 987 -1751
rect 896 -1817 909 -1753
rect 973 -1817 987 -1753
rect 1493 -1811 1506 -1747
rect 1570 -1811 1584 -1747
rect 1493 -1812 1584 -1811
rect 896 -1818 987 -1817
rect 900 -1820 980 -1818
rect 1500 -1820 1580 -1812
rect -820 -2443 -740 -2430
rect -820 -2499 -810 -2443
rect -754 -2499 -740 -2443
rect -820 -2510 -740 -2499
<< via3 >>
rect 1530 -457 1594 -453
rect 926 -550 990 -486
rect 1530 -513 1534 -457
rect 1534 -513 1590 -457
rect 1590 -513 1594 -457
rect 1530 -517 1594 -513
rect -287 -691 -223 -687
rect -287 -747 -283 -691
rect -283 -747 -227 -691
rect -227 -747 -223 -691
rect -287 -751 -223 -747
rect 312 -696 376 -692
rect 312 -752 316 -696
rect 316 -752 372 -696
rect 372 -752 376 -696
rect 312 -756 376 -752
rect 1561 -752 1625 -688
rect 2109 -694 2173 -690
rect 2109 -750 2113 -694
rect 2113 -750 2169 -694
rect 2169 -750 2173 -694
rect 2109 -754 2173 -750
rect 2710 -694 2774 -690
rect 2710 -750 2714 -694
rect 2714 -750 2770 -694
rect 2770 -750 2774 -694
rect 2710 -754 2774 -750
rect -292 -1119 -228 -1115
rect -292 -1175 -288 -1119
rect -288 -1175 -232 -1119
rect -232 -1175 -228 -1119
rect -292 -1179 -228 -1175
rect 278 -1112 342 -1106
rect 278 -1168 283 -1112
rect 283 -1168 339 -1112
rect 339 -1168 342 -1112
rect 278 -1170 342 -1168
rect 906 -1114 970 -1110
rect 906 -1170 910 -1114
rect 910 -1170 966 -1114
rect 966 -1170 970 -1114
rect 906 -1174 970 -1170
rect -288 -1538 -224 -1534
rect -288 -1594 -284 -1538
rect -284 -1594 -228 -1538
rect -228 -1594 -224 -1538
rect -288 -1598 -224 -1594
rect 281 -1534 345 -1528
rect 281 -1590 284 -1534
rect 284 -1590 340 -1534
rect 340 -1590 345 -1534
rect 281 -1592 345 -1590
rect 2111 -1112 2175 -1108
rect 2111 -1168 2115 -1112
rect 2115 -1168 2171 -1112
rect 2171 -1168 2175 -1112
rect 2111 -1172 2175 -1168
rect 2711 -1111 2775 -1107
rect 2711 -1167 2715 -1111
rect 2715 -1167 2771 -1111
rect 2771 -1167 2775 -1111
rect 2711 -1171 2775 -1167
rect 1222 -1284 1286 -1280
rect 1222 -1340 1226 -1284
rect 1226 -1340 1282 -1284
rect 1282 -1340 1286 -1284
rect 1222 -1344 1286 -1340
rect 3386 -1333 3450 -1329
rect 3386 -1389 3390 -1333
rect 3390 -1389 3446 -1333
rect 3446 -1389 3450 -1333
rect 3386 -1393 3450 -1389
rect 2105 -1542 2169 -1538
rect 2105 -1598 2109 -1542
rect 2109 -1598 2165 -1542
rect 2165 -1598 2169 -1542
rect 2105 -1602 2169 -1598
rect 2715 -1537 2779 -1533
rect 2715 -1593 2719 -1537
rect 2719 -1593 2775 -1537
rect 2775 -1593 2779 -1537
rect 2715 -1597 2779 -1593
rect 909 -1817 973 -1753
rect 1506 -1811 1570 -1747
<< metal4 >>
rect 1500 -453 1640 -440
rect 1500 -480 1530 -453
rect 900 -486 1530 -480
rect 900 -550 926 -486
rect 990 -517 1530 -486
rect 1594 -517 1640 -453
rect 990 -550 1640 -517
rect 900 -560 1640 -550
rect -289 -680 -221 -677
rect 906 -680 974 -666
rect 1559 -680 1627 -678
rect -1600 -687 3160 -680
rect -1600 -751 -287 -687
rect -223 -688 3160 -687
rect -223 -692 1561 -688
rect -223 -751 312 -692
rect -1600 -756 312 -751
rect 376 -752 1561 -692
rect 1625 -690 3160 -688
rect 1625 -752 2109 -690
rect 376 -754 2109 -752
rect 2173 -754 2710 -690
rect 2774 -754 3160 -690
rect 376 -756 3160 -754
rect -1600 -760 3160 -756
rect 310 -765 378 -760
rect 1559 -761 1627 -760
rect 2107 -763 2175 -760
rect 2708 -763 2776 -760
rect 276 -1100 344 -1096
rect 2109 -1100 2177 -1098
rect 2709 -1100 2777 -1097
rect -1600 -1106 3160 -1100
rect -1600 -1115 278 -1106
rect -1600 -1179 -292 -1115
rect -228 -1170 278 -1115
rect 342 -1107 3160 -1106
rect 342 -1108 2711 -1107
rect 342 -1110 2111 -1108
rect 342 -1170 906 -1110
rect -228 -1174 906 -1170
rect 970 -1172 2111 -1110
rect 2175 -1171 2711 -1108
rect 2775 -1171 3160 -1107
rect 2175 -1172 3160 -1171
rect 970 -1174 3160 -1172
rect -228 -1179 3160 -1174
rect -1600 -1180 3160 -1179
rect -294 -1188 -226 -1180
rect 904 -1183 972 -1180
rect 2109 -1181 2177 -1180
rect 1060 -1280 1459 -1246
rect 1060 -1324 1222 -1280
rect 1055 -1344 1222 -1324
rect 1286 -1324 1459 -1280
rect 3384 -1324 3452 -1319
rect 1286 -1329 3459 -1324
rect 1286 -1344 3386 -1329
rect 1055 -1393 3386 -1344
rect 3450 -1393 3459 -1329
rect 1055 -1401 3459 -1393
rect 3384 -1402 3452 -1401
rect 279 -1520 347 -1518
rect -1600 -1528 3160 -1520
rect -1600 -1534 281 -1528
rect -1600 -1598 -288 -1534
rect -224 -1592 281 -1534
rect 345 -1533 3160 -1528
rect 345 -1538 2715 -1533
rect 345 -1592 2105 -1538
rect -224 -1598 2105 -1592
rect -1600 -1600 2105 -1598
rect -290 -1607 -222 -1600
rect 279 -1601 347 -1600
rect 2103 -1602 2105 -1600
rect 2169 -1597 2715 -1538
rect 2779 -1597 3160 -1533
rect 2169 -1600 3160 -1597
rect 2169 -1602 2171 -1600
rect 2103 -1611 2171 -1602
rect 2713 -1606 2781 -1600
rect 900 -1747 1580 -1740
rect 900 -1753 1506 -1747
rect 900 -1817 909 -1753
rect 973 -1811 1506 -1753
rect 1570 -1811 1580 -1747
rect 973 -1817 1580 -1811
rect 900 -1820 1580 -1817
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_0
timestamp 1757161594
transform 0 1 -502 -1 0 -306
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_1
timestamp 1757161594
transform 0 1 -502 -1 0 -726
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_2
timestamp 1757161594
transform 0 1 698 -1 0 -726
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_3
timestamp 1757161594
transform 0 1 1898 -1 0 -726
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_4
timestamp 1757161594
transform 0 1 1298 -1 0 -726
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_5
timestamp 1757161594
transform 0 1 2498 -1 0 -726
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_6
timestamp 1757161594
transform 0 1 2498 -1 0 -306
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_7
timestamp 1757161594
transform 0 1 1898 -1 0 -306
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_8
timestamp 1757161594
transform 0 1 1298 -1 0 -306
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_9
timestamp 1757161594
transform 0 1 698 -1 0 -306
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_10
timestamp 1757161594
transform 0 1 98 -1 0 -306
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_11
timestamp 1757161594
transform 0 1 98 -1 0 -726
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_12
timestamp 1757161594
transform 0 1 1298 -1 0 -1566
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_13
timestamp 1757161594
transform 0 1 -502 -1 0 -1146
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_14
timestamp 1757161594
transform 0 1 98 -1 0 -1146
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_15
timestamp 1757161594
transform 0 1 698 -1 0 -1146
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_16
timestamp 1757161594
transform 0 1 1298 -1 0 -1146
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_17
timestamp 1757161594
transform 0 1 1898 -1 0 -1146
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_18
timestamp 1757161594
transform 0 1 2498 -1 0 -1146
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_19
timestamp 1757161594
transform 0 1 -502 -1 0 -1566
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_20
timestamp 1757161594
transform 0 1 98 -1 0 -1566
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_21
timestamp 1757161594
transform 0 1 698 -1 0 -1566
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_22
timestamp 1757161594
transform 0 1 98 -1 0 -1986
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_23
timestamp 1757161594
transform 0 1 1898 -1 0 -1566
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_24
timestamp 1757161594
transform 0 1 2498 -1 0 -1566
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_26
timestamp 1757161594
transform 0 1 1298 -1 0 -1986
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_27
timestamp 1757161594
transform 0 1 698 -1 0 -1986
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_28
timestamp 1757161594
transform 0 1 2498 -1 0 -1986
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_29
timestamp 1757161594
transform 0 1 1898 -1 0 -1986
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J88B3D  sky130_fd_pr__pfet_01v8_lvt_J88B3D_30
timestamp 1757161594
transform 0 1 -502 -1 0 -1986
box -194 -298 194 264
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_0
timestamp 1757161594
transform 0 1 -1002 -1 0 -1986
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_1
timestamp 1757161594
transform 0 1 -1002 -1 0 -1566
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_2
timestamp 1757161594
transform 0 1 -1002 -1 0 -1126
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_3
timestamp 1757161594
transform 0 1 -1002 -1 0 -706
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_4
timestamp 1757161594
transform 0 1 2998 -1 0 -1986
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_5
timestamp 1757161594
transform 0 1 -1002 -1 0 -306
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_6
timestamp 1757161594
transform 0 1 2998 -1 0 -1566
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_7
timestamp 1757161594
transform 0 1 2998 -1 0 -1146
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_8
timestamp 1757161594
transform 0 1 2998 -1 0 -726
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_9
timestamp 1757161594
transform 0 1 2998 -1 0 -306
box -194 -198 194 164
<< end >>
