* NGSPICE file created from op_amp_lvs_final.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_lvt_MTZNSY a_50_n136# a_n108_n136# a_n50_n162# w_n144_n198#
X0 a_50_n136# a_n50_n162# a_n108_n136# w_n144_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_KVZN99 w_n594_n198# a_500_n136# a_n558_n136# a_n500_n162#
X0 a_500_n136# a_n500_n162# a_n558_n136# w_n594_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
.ends

.subckt cs_p_5 w_n153_n413# m1_170_n270# m1_1670_4650# Vb
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_5 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_0 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_6 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_10 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_21 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_32 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_43 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_54 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_76 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_65 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_10 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_1 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_7 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_11 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_22 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_33 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_44 w_n153_n413# m1_170_n270# m1_1670_4650# Vb
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_55 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_77 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_66 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_11 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_2 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_12 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_23 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_34 w_n153_n413# m1_170_n270# m1_1670_4650# Vb
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_45 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_56 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_78 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_67 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_8 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_3 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_12 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_9 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_13 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_24 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_35 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_46 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_57 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_79 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_68 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_13 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_4 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_14 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_25 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_36 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_47 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_58 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_69 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_5 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_14 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_15 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_26 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_37 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_48 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_59 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_15 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_6 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_16 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_27 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_38 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_49 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_16 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_7 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_17 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_28 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_39 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_17 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_8 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_18 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_29 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_18 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_9 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_19 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_19 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_0 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_70 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_71 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_60 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_1 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_2 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_50 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_72 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_61 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_40 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_51 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_73 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_62 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_3 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_MTZNSY_4 m1_170_n270# m1_170_n270# m1_170_n270# w_n153_n413#
+ sky130_fd_pr__pfet_01v8_lvt_MTZNSY
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_30 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_41 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_52 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_74 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_63 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_20 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_31 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_42 w_n153_n413# m1_170_n270# m1_170_n270# m1_170_n270#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_53 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_75 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_64 w_n153_n413# m1_170_n270# Vb Vb sky130_fd_pr__pfet_01v8_lvt_KVZN99
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_BX6RT7 a_n108_n81# a_50_n81# a_n50_n107# VSUBS
X0 a_50_n81# a_n50_n107# a_n108_n81# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_N42WW9 a_n2000_n107# a_2000_n81# a_n2058_n81#
+ VSUBS
X0 a_2000_n81# a_n2000_n107# a_n2058_n81# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=20
.ends

.subckt block03 sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS m1_n144_4165# m1_n288_4065#
+ m1_n580_n270#
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_10 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_11 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_0 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_1 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_N42WW9_1 m1_n144_4165# m1_n580_n270# m1_n144_4165# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_N42WW9
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_2 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_N42WW9_0 m1_n144_4165# m1_n580_n270# m1_n288_4065# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_N42WW9
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_4 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_N42WW9_2 m1_n144_4165# m1_n580_n270# m1_n144_4165# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_N42WW9
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_3 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_N42WW9_3 m1_n144_4165# m1_n580_n270# m1_n288_4065# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_N42WW9
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_5 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_N42WW9_4 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_N42WW9
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_6 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_7 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_N42WW9_5 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_N42WW9
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_8 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
Xsky130_fd_pr__nfet_01v8_lvt_BX6RT7_9 m1_n580_n270# m1_n580_n270# m1_n580_n270# sky130_fd_pr__nfet_01v8_lvt_N42WW9_5/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_BX6RT7
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_J88B3D a_100_n236# a_n158_n236# a_n100_n262# w_n194_n298#
X0 a_100_n236# a_n100_n262# a_n158_n236# w_n194_n298# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_J8833D w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt block01 m1_n299_n1606# m1_n298_n759# m1_n595_n1313# m1_n303_n1187# m1_n581_n1736#
+ w_n1380_n2320#
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_0 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_1 m1_n581_n1736# w_n1380_n2320# m1_n298_n759#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_2 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_3 m1_n581_n1736# w_n1380_n2320# m1_n298_n759#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_4 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_5 m1_n581_n1736# w_n1380_n2320# m1_n298_n759#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_6 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_7 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_8 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_9 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_30 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_20 m1_n581_n1736# w_n1380_n2320# m1_n299_n1606#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_10 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_21 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_11 m1_n581_n1736# w_n1380_n2320# m1_n298_n759#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_22 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_23 m1_n581_n1736# w_n1380_n2320# m1_n299_n1606#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_12 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_14 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_13 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_24 m1_n581_n1736# w_n1380_n2320# m1_n299_n1606#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_15 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_26 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_16 m1_n581_n1736# w_n1380_n2320# m1_n298_n759#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_27 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_17 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_28 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_18 m1_n595_n1313# w_n1380_n2320# m1_n303_n1187#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_29 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J88B3D_19 m1_n581_n1736# w_n1380_n2320# m1_n299_n1606#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J88B3D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_0 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_1 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_3 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_2 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_4 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_5 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_6 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_7 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_8 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_9 w_n1380_n2320# w_n1380_n2320# w_n1380_n2320#
+ w_n1380_n2320# sky130_fd_pr__pfet_01v8_lvt_J8833D
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_LTPL8U a_n100_n117# a_100_n91# a_n158_n91# VSUBS
X0 a_100_n91# a_n100_n117# a_n158_n91# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.174 pd=1.78 as=0.174 ps=1.78 w=0.6 l=1
.ends

.subckt nmos_08 m1_450_510# m1_310_690# m1_0_0# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_0 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_1 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_2 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_3 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_5 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_4 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_6 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_7 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_10 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_8 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_11 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_12 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_9 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_13 m1_450_510# m1_310_690# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_14 m1_450_510# m1_450_510# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_15 m1_450_510# m1_450_510# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_17 m1_0_0# m1_0_0# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
Xsky130_fd_pr__nfet_01v8_lvt_LTPL8U_16 m1_450_510# m1_310_690# m1_0_0# VSUBS sky130_fd_pr__nfet_01v8_lvt_LTPL8U
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_34DASA a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt block02 m1_n552_n4379# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530#
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_10 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_21 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_32 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_11 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_22 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_33 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_12 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_23 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_34 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_13 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_24 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_35 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_14 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_36 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_25 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_16 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_15 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_37 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_38 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_27 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_26 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_0 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS m1_n350_n4530#
+ m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_17 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_39 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_28 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_1 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_18 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_29 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_2 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_19 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_4 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_3 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_5 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_6 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_7 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_8 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_9 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_30 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n552_n4379# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_20 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ m1_n350_n4530# m1_n560_n3972# sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
Xsky130_fd_pr__nfet_01v8_lvt_34DASA_31 sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_34DASA_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_34DASA
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_MYAC2F m3_n1186_n540# c1_n1146_n500#
X0 c1_n1146_n500# m3_n1186_n540# sky130_fd_pr__cap_mim_m3_1 l=5 w=10
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_DP2CMY c1_n646_n1000# m3_n686_n1040#
X0 c1_n646_n1000# m3_n686_n1040# sky130_fd_pr__cap_mim_m3_1 l=10 w=5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_G6WD7P m3_n686_n540# c1_n646_n500#
X0 c1_n646_n500# m3_n686_n540# sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_GQMTM9 m3_n1186_n1040# c1_n1146_n1000#
X0 c1_n1146_n1000# m3_n1186_n1040# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_B9M9HY m3_n1186_n1040# c1_n1146_n1000#
X0 c1_n1146_n1000# m3_n1186_n1040# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
.ends

.subckt cap m4_6650_4870# m4_8770_5032# m4_8940_7520# m4_6540_2680# m4_9320_1970#
Xsky130_fd_pr__cap_mim_m3_1_MYAC2F_2 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_MYAC2F
Xsky130_fd_pr__cap_mim_m3_1_MYAC2F_3 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_MYAC2F
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_0 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_2 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_1 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_3 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_4 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_5 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_6 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_G6WD7P_0 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_G6WD7P
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_7 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_G6WD7P_1 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_G6WD7P
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_8 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_G6WD7P_2 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_G6WD7P
Xsky130_fd_pr__cap_mim_m3_1_G6WD7P_3 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_G6WD7P
Xsky130_fd_pr__cap_mim_m3_1_DP2CMY_9 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_DP2CMY
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_15 m4_8940_7520# m4_8770_5032# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_1 m4_8940_7520# m4_8770_5032# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_17 m4_8940_7520# m4_8770_5032# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_3 m4_6650_4870# m4_6540_2680# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_18 m4_6650_4870# m4_6540_2680# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_4 m4_6650_4870# m4_6540_2680# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_19 m4_6650_4870# m4_6540_2680# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_B9M9HY_0 m4_8940_7520# m4_8770_5032# sky130_fd_pr__cap_mim_m3_1_B9M9HY
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_5 m4_6650_4870# m4_6540_2680# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_GQMTM9_6 m4_8940_7520# m4_8770_5032# sky130_fd_pr__cap_mim_m3_1_GQMTM9
Xsky130_fd_pr__cap_mim_m3_1_MYAC2F_0 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_MYAC2F
Xsky130_fd_pr__cap_mim_m3_1_MYAC2F_1 m4_9320_1970# m4_9320_1970# sky130_fd_pr__cap_mim_m3_1_MYAC2F
.ends

.subckt sky130_fd_pr__res_generic_po_RETGBZ a_n50_n4430# a_n50_4000#
X0 a_n50_4000# a_n50_n4430# sky130_fd_pr__res_generic_po w=0.5 l=40
.ends

.subckt res m1_10_8850# m1_160_8700# m1_5710_8850#
Xsky130_fd_pr__res_generic_po_RETGBZ_40 m1_5560_0# m1_5710_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_30 m1_3010_n110# m1_3310_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_0 m1_1960_0# m1_2260_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_32 m1_4810_n110# m1_4510_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_21 m1_4360_0# m1_4060_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_20 m1_4210_n110# m1_3910_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_31 m1_3160_0# m1_3460_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_1 m1_1810_n110# m1_1510_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_10 m1_610_n110# m1_910_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_33 m1_4960_0# m1_4660_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_22 m1_4210_n110# m1_4510_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_2 m1_1960_0# m1_1660_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_11 m1_760_0# m1_1060_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_34 m1_4810_n110# m1_5110_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_23 m1_4360_0# m1_4660_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_3 m1_1810_n110# m1_2110_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_12 m1_160_0# m1_460_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_35 m1_4960_0# m1_5260_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_24 m1_2410_n110# m1_2110_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_4 m1_1360_0# m1_1660_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_13 m1_10_n110# m1_310_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_36 m1_5410_n110# m1_5110_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_25 m1_2560_0# m1_2260_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_5 m1_1210_n110# m1_1510_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_14 m1_160_0# m1_160_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_37 m1_5560_0# m1_5260_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_26 m1_2410_n110# m1_2710_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_6 m1_1360_0# m1_1060_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_15 m1_10_n110# m1_10_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_38 m1_5410_n110# m1_5710_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_16 m1_3610_n110# m1_3310_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_27 m1_2560_0# m1_2860_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_7 m1_1210_n110# m1_910_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_18 m1_3610_n110# m1_3910_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_17 m1_3760_0# m1_3460_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_29 m1_3160_0# m1_2860_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_28 m1_3010_n110# m1_2710_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_9 m1_760_0# m1_460_8700# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_8 m1_610_n110# m1_310_8850# sky130_fd_pr__res_generic_po_RETGBZ
Xsky130_fd_pr__res_generic_po_RETGBZ_19 m1_3760_0# m1_4060_8700# sky130_fd_pr__res_generic_po_RETGBZ
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_LHHU6U a_n108_n86# w_n144_n148# a_50_n86# a_n50_n112#
X0 a_50_n86# a_n50_n112# a_n108_n86# w_n144_n148# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_W2HEQA a_n1000_n112# a_1000_n86# a_n1058_n86#
+ w_n1094_n148#
X0 a_1000_n86# a_n1000_n112# a_n1058_n86# w_n1094_n148# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=10
.ends

.subckt block04 m1_193_n116# m1_51_n253# m1_n570_220# m1_598_4# m1_n450_n2340# m1_456_124#
+ w_n500_n2860#
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_6 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_7 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_8 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_9 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_10 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_11 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_10 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_11 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_0 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_1 m1_193_n116# m1_n450_n2340# m1_51_n253# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_2 m1_598_4# m1_456_124# m1_51_n253# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_3 m1_598_4# m1_456_124# m1_51_n253# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_4 m1_193_n116# m1_n450_n2340# m1_51_n253# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_5 m1_193_n116# m1_n450_n2340# m1_51_n253# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_6 m1_598_4# m1_456_124# m1_51_n253# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_8 m1_193_n116# m1_n450_n2340# m1_51_n253# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_7 m1_598_4# m1_456_124# m1_51_n253# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_W2HEQA_9 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_W2HEQA
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_0 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_2 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_1 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_3 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_4 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
Xsky130_fd_pr__pfet_01v8_lvt_LHHU6U_5 w_n500_n2860# w_n500_n2860# w_n500_n2860# w_n500_n2860#
+ sky130_fd_pr__pfet_01v8_lvt_LHHU6U
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_6DE3T6 a_15_n131# a_n33_91# a_n73_n131# VSUBS
X0 a_15_n131# a_n33_91# a_n73_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt switchblock beta Vbias1 Vbias2 Vbias3 Vbias4 en_1 en_2 m1_n330_n2520# m1_140_n2620#
+ m1_n330_n2220# m1_140_n2020# sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS w_n12993_n4583#
+ m1_n330_n720# m1_n330_n120# m1_n330_n1320# m1_140_n1420# m1_140_n820# m1_140_n220#
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_0 m1_140_n2620# en_2 m1_n330_n2520# sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_1 m1_140_n2620# en_1 beta sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_2 m1_140_n2020# en_1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_3 m1_140_n2020# en_2 m1_n330_n2220# sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_4 m1_140_n1420# en_1 Vbias2 sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_5 m1_140_n820# en_1 Vbias3 sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_6 m1_140_n1420# en_2 m1_n330_n1320# sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_7 m1_140_n220# en_1 Vbias4 sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_8 m1_140_n820# en_2 m1_n330_n720# sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
Xsky130_fd_pr__nfet_01v8_lvt_6DE3T6_9 m1_140_n220# en_2 m1_n330_n120# sky130_fd_pr__nfet_01v8_lvt_6DE3T6_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_6DE3T6
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_U8838H a_100_n536# a_n158_n536# a_n100_n562# w_n194_n598#
X0 a_100_n536# a_n100_n562# a_n158_n536# w_n194_n598# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=1
.ends

.subckt switchblock01 w_n480_n1940# m1_820_n900# m1_1320_n900# m1_n390_n60# m1_n270_n180#
+ m1_n150_n300#
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_10 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_10 m1_820_n900# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_11 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_11 m1_n390_n60# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_12 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_12 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_13 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_13 m1_n150_n300# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_0 m1_1320_n900# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_14 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_15 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_1 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_14 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_2 m1_n270_n180# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_15 m1_n270_n180# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_3 m1_n390_n60# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_4 m1_n150_n300# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_5 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_7 m1_820_n900# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_6 m1_1320_n900# w_n480_n1940# m1_n150_n300# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_8 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_U8838H_9 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_U8838H
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_0 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_1 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_2 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_3 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_4 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_5 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_6 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_7 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_8 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
Xsky130_fd_pr__pfet_01v8_lvt_J8833D_9 w_n480_n1940# w_n480_n1940# w_n480_n1940# w_n480_n1940#
+ sky130_fd_pr__pfet_01v8_lvt_J8833D
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_NVX44G a_200_n536# w_n396_n684# a_n258_n536# a_n200_n562#
+ li_n360_n648#
X0 a_200_n536# a_n200_n562# a_n258_n536# w_n396_n684# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_LVXMRT a_n2000_n161# w_n2196_n284# a_2000_n64#
+ a_n2058_n64#
X0 a_2000_n64# a_n2000_n161# a_n2058_n64# w_n2196_n284# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ZVWESF a_200_n531# a_n200_n557# a_n258_n531# a_n360_n643#
+ li_n360_n643#
X0 a_200_n531# a_n200_n557# a_n258_n531# a_n360_n643# sky130_fd_pr__nfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_2QSR6E a_200_n236# w_n396_n384# a_n258_n236# a_n200_n262#
X0 a_200_n236# a_n200_n262# a_n258_n236# w_n396_n384# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_JY4D7E a_200_n236# w_n396_n384# a_n258_n236# a_n200_n262#
+ li_n360_n348#
X0 a_200_n236# a_n200_n262# a_n258_n236# w_n396_n384# sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_VYCASF a_200_n231# a_n200_n257# a_n258_n231# a_n360_n343#
+ li_n360_n343#
X0 a_200_n231# a_n200_n257# a_n258_n231# a_n360_n343# sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_V2BN2G a_200_n231# a_n200_n257# a_n258_n231# a_n360_n343#
X0 a_200_n231# a_n200_n257# a_n258_n231# a_n360_n343# sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_UY454G a_200_n536# w_n396_n684# a_n258_n536# a_n200_n562#
+ li_n360_n648#
X0 a_200_n536# a_n200_n562# a_n258_n536# w_n396_n684# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.58 as=1.45 ps=10.58 w=5 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_9UXMRD a_n2000_n161# li_n2160_n248# w_n2196_n284#
+ a_2000_n64# a_n2058_n64#
X0 a_2000_n64# a_n2000_n161# a_n2058_n64# w_n2196_n284# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_PAU7SL a_100_n169# a_n260_n343# a_n158_n169# a_n100_n257#
X0 a_100_n169# a_n100_n257# a_n158_n169# a_n260_n343# sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt bias_dummy Vbias1 Vbias2 Vbias3 Vbias4 m1_3751_n8170# M46_4/VSUBS a_2860_n8920#
+ PBias w_1870_n4070#
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_6 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM43_1 Vbias1 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM42_B m1_1890_n4940# w_1870_n4070# m1_1890_n4940# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_LVXMRT
XM35_A m1_3751_n8170# m1_2980_n7670# m1_2980_n7670# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_7 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM43_2 Vbias1 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM35_B m1_3751_n8170# m1_2980_n7670# m1_2980_n7670# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_8 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM43_3 Vbias1 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM35_C m1_3751_n8170# m1_2980_n7670# m1_2980_n7670# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_9 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM43_4 Vbias1 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM33_A M46_4/VSUBS m1_2100_n5010# m1_2100_n5010# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
XM35_D m1_3751_n8170# m1_2980_n7670# m1_2980_n7670# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__pfet_01v8_lvt_2QSR6E_0 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ sky130_fd_pr__pfet_01v8_lvt_2QSR6E
XM35_E m1_3751_n8170# m1_2980_n7670# m1_2980_n7670# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_0 m1_3751_n8170# m1_2980_n7670# m1_2980_n7670#
+ M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
XM33_B M46_4/VSUBS m1_2100_n5010# m1_2100_n5010# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
XM35_F m1_3751_n8170# m1_2980_n7670# m1_2980_n7670# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_1 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
XM35_G m1_3751_n8170# m1_2980_n7670# m1_2980_n7670# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_2 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_3 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_4 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_5 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_6 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_0 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_7 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_1 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
Xsky130_fd_pr__nfet_01v8_lvt_ZVWESF_8 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_2 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
XM38_A PBias w_1870_n4070# w_1870_n4070# m1_2870_n6990# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_10 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
XM46_2 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_3 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
XM38_B PBias w_1870_n4070# w_1870_n4070# m1_2870_n6990# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_11 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
XM46_3 Vbias4 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM38_C PBias w_1870_n4070# w_1870_n4070# m1_2870_n6990# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM44_1 Vbias2 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM46_4 Vbias4 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_5 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
XM36_A M46_4/VSUBS m1_2980_n7670# m1_2870_n6990# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
XM38_D PBias w_1870_n4070# w_1870_n4070# m1_2870_n6990# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_6 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
XM44_2 Vbias2 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM36_B M46_4/VSUBS m1_2980_n7670# m1_2870_n6990# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
XM44_3 Vbias2 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_7 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
XM41_A M46_4/VSUBS m1_2100_n5010# m1_1890_n4940# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_8 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
XM44_4 Vbias2 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM41_B M46_4/VSUBS m1_2100_n5010# m1_1890_n4940# M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
XM34_A m1_2980_n7670# w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_9 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
XM34_B m1_2980_n7670# w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM34_C m1_2980_n7670# w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM34_D m1_2980_n7670# w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_10 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM32_A m1_2100_n5010# w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_11 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_V2BN2G_0 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_V2BN2G
XM32_B m1_2100_n5010# w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_12 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM32_C m1_2100_n5010# w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_0 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_13 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM32_D m1_2100_n5010# w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_1 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_14 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_2 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
Xsky130_fd_pr__pfet_01v8_lvt_UY454G_0 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_UY454G
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_15 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_3 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_16 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_4 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_0 Vbias4 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070#
+ sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM39_A m1_2870_n6990# w_1870_n4070# w_1870_n4070# m1_2870_n6990# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_5 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_1 Vbias4 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070#
+ sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM39_B m1_2870_n6990# w_1870_n4070# w_1870_n4070# m1_2870_n6990# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM39_C m1_2870_n6990# w_1870_n4070# w_1870_n4070# m1_2870_n6990# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_7 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_3 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM45_1 Vbias3 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM39_D m1_2870_n6990# w_1870_n4070# w_1870_n4070# m1_2870_n6990# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_8 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
XM37_A M46_4/VSUBS m1_2100_n5010# PBias M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
XM45_2 Vbias3 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_10 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_4 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM37_B M46_4/VSUBS m1_2100_n5010# PBias M46_4/VSUBS M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_ZVWESF
Xsky130_fd_pr__nfet_01v8_lvt_VYCASF_9 M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS M46_4/VSUBS
+ M46_4/VSUBS sky130_fd_pr__nfet_01v8_lvt_VYCASF
Xsky130_fd_pr__pfet_01v8_lvt_NVX44G_5 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
XM45_3 Vbias3 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
Xsky130_fd_pr__pfet_01v8_lvt_JY4D7E_11 w_1870_n4070# w_1870_n4070# w_1870_n4070# w_1870_n4070#
+ w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_JY4D7E
XM42_A m1_1890_n4940# w_1870_n4070# w_1870_n4070# m1_1890_n4940# w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_9UXMRD
XM40 m1_2100_n5010# M46_4/VSUBS PBias m1_1890_n4940# sky130_fd_pr__nfet_01v8_lvt_PAU7SL
XM45_4 Vbias3 w_1870_n4070# w_1870_n4070# PBias w_1870_n4070# sky130_fd_pr__pfet_01v8_lvt_NVX44G
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_VVFJJL a_n1000_n257# a_1000_n231# a_n1058_n231#
+ VSUBS
X0 a_1000_n231# a_n1000_n257# a_n1058_n231# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_ND6TEZ a_n158_n231# a_100_n231# a_n100_n257# VSUBS
X0 a_100_n231# a_n100_n257# a_n158_n231# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt diff_in_03 m1_70_0# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS a_1820_4690#
+ m1_40_4430# m1_n100_n530# in- in+
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_18 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_19 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_7 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_8 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_9 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_20 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_21 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_10 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_22 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_11 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_12 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_14 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_13 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_25 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_24 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_15 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_16 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_17 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_0 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_18 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_19 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_2 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_3 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_5 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_4 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_6 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_10 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_20 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_21 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_7 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_22 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_8 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_12 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_0 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_ND6TEZ_9 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_ND6TEZ
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_1 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_13 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_2 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_24 a_1820_4690# a_1820_4690# a_1820_4690# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_14 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_25 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_3 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_15 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_4 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_16 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_5 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_17 in+ m1_70_0# m1_n100_n530# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
Xsky130_fd_pr__nfet_01v8_lvt_VVFJJL_6 in- m1_70_0# m1_40_4430# sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_VVFJJL
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_76U4T2 a_1000_n136# w_n1094_n198# a_n1058_n136#
+ a_n1000_n162#
X0 a_1000_n136# a_n1000_n162# a_n1058_n136# w_n1094_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_KVZWZ9 w_n194_n198# a_100_n136# a_n158_n136# a_n100_n162#
X0 a_100_n136# a_n100_n162# a_n158_n136# w_n194_n198# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt pmos_07 m1_730_40# m1_480_40# w_n80_n500# m1_100_n80#
Xsky130_fd_pr__pfet_01v8_lvt_76U4T2_0 m1_100_n80# w_n80_n500# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_76U4T2
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_10 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_76U4T2_1 m1_480_40# w_n80_n500# m1_100_n80# m1_730_40#
+ sky130_fd_pr__pfet_01v8_lvt_76U4T2
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_11 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_76U4T2_2 m1_480_40# w_n80_n500# m1_100_n80# m1_730_40#
+ sky130_fd_pr__pfet_01v8_lvt_76U4T2
Xsky130_fd_pr__pfet_01v8_lvt_76U4T2_4 m1_730_40# w_n80_n500# m1_100_n80# m1_730_40#
+ sky130_fd_pr__pfet_01v8_lvt_76U4T2
Xsky130_fd_pr__pfet_01v8_lvt_76U4T2_5 m1_730_40# w_n80_n500# m1_100_n80# m1_730_40#
+ sky130_fd_pr__pfet_01v8_lvt_76U4T2
Xsky130_fd_pr__pfet_01v8_lvt_76U4T2_6 m1_100_n80# w_n80_n500# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_76U4T2
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_0 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_1 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_2 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_3 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_4 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_5 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_6 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_7 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_9 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_8 w_n80_n500# m1_100_n80# m1_100_n80# m1_100_n80#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_RSMGKB a_n108_n86# w_n144_n148# a_50_n86# a_n50_n112#
X0 a_50_n86# a_n50_n112# a_n108_n86# w_n144_n148# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_RSW4TG a_n1000_n112# a_1000_n86# a_n1058_n86#
+ w_n1094_n148#
X0 a_1000_n86# a_n1000_n112# a_n1058_n86# w_n1094_n148# sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=10
.ends

.subckt pmos_05 m1_n70_2090# w_6467_5190# w_6447_n690# m1_360_2270# w_n313_n573# w_6697_n690#
+ m1_360_40# m1_370_4410# w_6707_5190# m1_57_5130# Vbin
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_16 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_9 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_38 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_7 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_17 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_39 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_28 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_8 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_18 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_9 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_29 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_19 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_60 m1_57_5130# m1_57_5130# m1_57_5130# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_61 m1_57_5130# m1_57_5130# m1_57_5130# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_62 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_50 Vbin m1_57_5130# Vbin w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_51 Vbin m1_57_5130# Vbin w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_63 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_52 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_64 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_53 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_20 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_65 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_54 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_21 m1_57_5130# m1_57_5130# m1_57_5130# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_10 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_55 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_44 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_22 m1_57_5130# m1_57_5130# m1_57_5130# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_11 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_56 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_45 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_12 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_23 m1_57_5130# m1_57_5130# m1_57_5130# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_57 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_46 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_13 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_58 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_47 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_14 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_59 Vbin m1_57_5130# Vbin w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_16 Vbin m1_57_5130# Vbin w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_15 m1_57_5130# m1_57_5130# m1_57_5130# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_17 Vbin m1_57_5130# Vbin w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_18 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_19 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_40 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_0 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_1 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_41 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_30 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_2 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_20 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_42 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_0 Vbin m1_57_5130# Vbin w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_31 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_3 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_21 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_10 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_43 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_32 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_1 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_4 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_11 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_22 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_44 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_33 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_2 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_5 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_12 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_6 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_23 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_34 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_3 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_13 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_14 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_7 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_24 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_25 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_36 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_35 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_4 Vbin m1_370_4410# m1_360_2270# w_n313_n573#
+ sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_15 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_8 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_26 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSMGKB_37 m1_57_5130# w_n313_n573# m1_57_5130# m1_57_5130#
+ sky130_fd_pr__pfet_01v8_lvt_RSMGKB
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_5 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
Xsky130_fd_pr__pfet_01v8_lvt_RSW4TG_6 Vbin m1_n70_2090# m1_360_40# w_n313_n573# sky130_fd_pr__pfet_01v8_lvt_RSW4TG
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_G235U9 a_1000_n81# a_n1058_n81# a_n1000_n107#
+ VSUBS
X0 a_1000_n81# a_n1000_n107# a_n1058_n81# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_QGYFYD a_n108_n81# a_50_n81# a_n50_n107# VSUBS
X0 a_50_n81# a_n50_n107# a_n108_n81# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt diff_in_04 m1_290_4320# m1_360_6670# m1_290_0# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ m1_290_4520# m1_290_2060# Vref m1_0_n280# m1_410_2610#
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_8 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_9 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_0 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_1 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_2 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_3 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_5 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_4 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_6 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_7 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_40 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_41 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_30 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_8 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_42 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_31 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_20 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_43 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_32 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_21 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_9 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_10 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_44 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_33 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_22 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_11 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_45 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_34 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_12 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_23 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_20 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_46 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_24 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_35 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_13 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_21 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_10 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_47 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_36 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_25 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_14 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_22 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_11 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_12 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_37 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_26 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_15 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_23 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_13 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_39 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_38 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_27 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_28 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_16 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_17 m1_290_4320# m1_290_4520# m1_360_6670# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_14 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_29 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_18 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_19 m1_290_4320# m1_290_0# m1_410_2610# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_15 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_0 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_16 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_1 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_17 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_18 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_2 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGYFYD_19 m1_0_n280# m1_0_n280# m1_0_n280# sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGYFYD
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_3 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_4 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_5 m1_290_2060# m1_290_4520# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_6 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_7 m1_290_2060# m1_290_0# Vref sky130_fd_pr__nfet_01v8_lvt_QGYFYD_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_G235U9
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_F22EEM a_n1000_n157# a_1000_n131# a_n1058_n131#
+ VSUBS
X0 a_1000_n131# a_n1000_n157# a_n1058_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_6WKBEZ a_100_n131# a_n100_n157# a_n158_n131# VSUBS
X0 a_100_n131# a_n100_n157# a_n158_n131# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt nmos_cl_02 m1_1500_5160# m1_n250_n4820# m1_n110_1640# m1_2320_n2290# m1_2320_n4350#
+ Vbias2 m1_2130_4710# m4_n590_n5050# Vss m1_420_n2290# m1_420_2070#
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_90 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_80 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_91 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_70 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_81 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_93 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_60 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_71 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_82 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_94 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_50 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_72 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_83 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_61 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_40 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_95 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_51 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_73 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_84 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_62 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_41 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_30 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_63 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_52 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_85 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_42 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_31 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_64 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_53 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_75 Vbias2 Vbias2 Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_86 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_20 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_43 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_32 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_65 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_54 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_76 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_87 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_10 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_21 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_44 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_33 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_66 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_55 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_77 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_88 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_22 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_40 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_45 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_34 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_67 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_56 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_78 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_89 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_23 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_12 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_35 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_24 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_68 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_57 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_46 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_79 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_13 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_41 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_30 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_0 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_42 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_31 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_36 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_1 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_58 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_20 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_47 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_69 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_14 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_25 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_0 Vbias2 Vbias2 Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_37 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_59 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_48 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_15 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_26 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_43 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_32 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_2 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_10 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_21 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_1 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_38 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_3 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_49 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_16 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_27 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_44 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_33 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_11 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_22 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_2 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_39 Vbias2 m1_420_n2290# m1_n250_n4820# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_17 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_45 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_34 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_23 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_4 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_12 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_3 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_29 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_5 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_18 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_35 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_24 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_13 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_4 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_19 Vbias2 m1_2320_n2290# m1_2320_n4350# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_36 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_25 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_6 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_14 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_5 Vbias2 m1_420_2070# m1_2130_4710# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_7 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_37 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_26 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_15 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_6 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_38 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_27 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_8 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_16 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_7 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_39 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_28 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_9 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_17 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_8 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_29 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_18 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
Xsky130_fd_pr__nfet_01v8_lvt_F22EEM_9 Vbias2 m1_420_2070# m1_n110_1640# Vss sky130_fd_pr__nfet_01v8_lvt_F22EEM
Xsky130_fd_pr__nfet_01v8_lvt_6WKBEZ_19 Vss Vss Vss Vss sky130_fd_pr__nfet_01v8_lvt_6WKBEZ
.ends

.subckt pmos_06 w_n290_n530# Vin m1_60_n390# m1_n60_40# m1_470_n50#
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_10 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_21 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_0 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_11 w_n290_n530# m1_60_n390# m1_n60_40# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_1 w_n290_n530# m1_60_n390# m1_n60_40# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_12 w_n290_n530# m1_60_n390# m1_n60_40# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_2 w_n290_n530# m1_60_n390# m1_470_n50# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_20 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_21 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_13 w_n290_n530# m1_60_n390# m1_470_n50# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_3 w_n290_n530# m1_60_n390# m1_470_n50# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_14 w_n290_n530# m1_60_n390# m1_470_n50# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_4 w_n290_n530# m1_60_n390# m1_470_n50# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_12 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_15 w_n290_n530# m1_60_n390# m1_470_n50# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_5 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_13 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_16 w_n290_n530# m1_60_n390# m1_470_n50# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_7 w_n290_n530# m1_60_n390# m1_n60_40# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_6 w_n290_n530# m1_60_n390# m1_n60_40# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_14 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_17 w_n290_n530# m1_60_n390# m1_n60_40# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_18 w_n290_n530# m1_60_n390# m1_n60_40# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_8 w_n290_n530# m1_60_n390# m1_n60_40# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_15 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZN99_9 w_n290_n530# m1_60_n390# m1_470_n50# Vin sky130_fd_pr__pfet_01v8_lvt_KVZN99
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_16 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_17 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_18 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_19 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_0 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_1 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_2 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_3 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_4 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_5 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_6 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_7 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_9 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
Xsky130_fd_pr__pfet_01v8_lvt_KVZWZ9_8 w_n290_n530# m1_60_n390# m1_60_n390# m1_60_n390#
+ sky130_fd_pr__pfet_01v8_lvt_KVZWZ9
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_QGGREF a_n108_n81# a_50_n81# a_n50_n107# VSUBS
X0 a_50_n81# a_n50_n107# a_n108_n81# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
.ends

.subckt nmos_cload_01 m1_n390_n2330# m1_n390_2140# m4_6030_n2460# m1_n480_n2830# Vbias1
+ m1_590_n180# m1_1890_2150# m1_n300_n2420# a_n370_n2650# sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_8 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS m1_n300_n2420#
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_9 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS Vbias1
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_0 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_40 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_41 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_30 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_2 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_3 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_42 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_31 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_20 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_4 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_43 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_33 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_32 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_22 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_21 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_11 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_10 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_44 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_5 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_34 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_23 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_12 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_6 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_35 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_24 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_40 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n390_2140# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_41 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n300_n2420# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_13 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_30 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_7 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_36 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_25 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_20 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_590_n180# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_42 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_31 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_1890_2150# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_14 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_37 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_26 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_21 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_590_n180# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_10 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n300_n2420# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_43 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_15 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_32 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n300_n2420# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_9 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_38 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_27 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_22 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_11 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_1890_2150# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_16 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_33 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_44 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_39 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_28 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_12 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_23 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_17 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_34 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n480_n2830# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_29 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_13 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_19 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_QGGREF_18 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_QGGREF
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_35 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_24 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n390_n2330# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_14 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_36 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_25 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n390_n2330# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_37 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_26 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_590_n180# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_17 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n390_n2330# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_16 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n480_n2830# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_38 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_39 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n390_2140# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_27 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_28 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_18 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_n390_n2330# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_29 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ m1_590_n180# Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_19 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS
+ Vbias1 Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_0 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS Vbias1
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS Vbias1
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_2 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS Vbias1
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_3 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS Vbias1
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_4 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS m1_n390_2140#
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_5 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS m1_n390_2140#
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_6 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS Vbias1
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
Xsky130_fd_pr__nfet_01v8_lvt_G235U9_7 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS Vbias1
+ Vbias1 sky130_fd_pr__nfet_01v8_lvt_QGGREF_9/VSUBS sky130_fd_pr__nfet_01v8_lvt_G235U9
.ends

.subckt Diff_opamp_ly Vbias3 Vbias2 m1_7390_12740# nmos_cload_01_1/Vbias1 m3_7390_13910#
+ m1_5550_12740# diff_in_04_0/Vref a_5590_12246# a_14260_10340# m1_930_12740# m1_4090_12740#
+ a_2690_12256# diff_in_03_0/in- a_1590_5786# m1_2650_12740# li_12480_21783# nmos_cload_01_1/a_n370_n2650#
+ m3_7630_14190# diff_in_03_0/in+ a_21110_n524# w_12480_21783# m3_12530_14200# m1_12460_17310#
+ a_19140_n514# pmos_07_0/VSUBS m1_10860_12520# w_367_15127#
Xdiff_in_03_0 m2_8270_9210# pmos_07_0/VSUBS pmos_07_0/VSUBS m3_n60_15150# m3_220_15330#
+ diff_in_03_0/in- diff_in_03_0/in+ diff_in_03
Xnmos_08_0 Vbias3 pmos_05_0/Vbin pmos_07_0/VSUBS pmos_07_0/VSUBS nmos_08
Xpmos_07_0 m3_10960_15920# pmos_06_0/Vin w_367_15127# w_367_15127# pmos_07
Xpmos_05_0 m3_n60_15150# w_367_15127# w_367_15127# m3_7630_14190# w_367_15127# w_367_15127#
+ m3_7390_13910# m3_220_15330# w_367_15127# w_367_15127# pmos_05_0/Vbin pmos_05
Xdiff_in_04_0 m3_10960_15920# m3_7630_14190# m3_7460_n660# pmos_07_0/VSUBS m3_7460_n10#
+ pmos_06_0/Vin diff_in_04_0/Vref pmos_07_0/VSUBS m3_7390_13910# diff_in_04
Xnmos_cl_02_1 pmos_07_0/VSUBS m3_7460_5410# m3_7460_210# m3_7390_13910# m3_7460_5210#
+ Vbias2 m3_7460_410# m3_7460_410# pmos_07_0/VSUBS m3_7630_14190# m2_8270_9210# nmos_cl_02
Xpmos_06_0 w_367_15127# pmos_06_0/Vin w_367_15127# m3_n60_15150# m3_220_15330# pmos_06
Xnmos_cload_01_1 m3_7460_410# m3_7460_5210# m3_7460_210# m3_7460_n660# nmos_cload_01_1/Vbias1
+ m3_7460_5410# m3_7460_n10# m3_7460_210# nmos_cload_01_1/a_n370_n2650# pmos_07_0/VSUBS
+ nmos_cload_01
.ends

.subckt x2stage_op_amp m1_14500_16280# Diff_opamp_ly_0/li_12480_21783# m3_n7330_11130#
+ m2_n6630_12060# switchblock_1/en_2 switchblock_1/en_1 w_12480_17180# bias_dummy_0/PBias
+ m1_15020_16390# Diff_opamp_ly_0/diff_in_03_0/in+ Diff_opamp_ly_0/w_12480_21783#
+ w_12480_17590# Diff_opamp_ly_0/diff_in_04_0/Vref Diff_opamp_ly_0/diff_in_03_0/in-
+ w_12790_18670# cap_1/VSUBS w_12670_17180# m2_n6620_11820# m4_30310_15630# w_n610_16180#
+ Diff_opamp_ly_0/nmos_cload_01_1/a_n370_n2650#
Xcs_p_5_0 w_n610_16180# w_n610_16180# m3_17920_18750# cs_p_5_0/Vb cs_p_5
Xblock03_0 cap_1/VSUBS m1_20390_14580# m1_20250_14460# cap_1/VSUBS block03
Xblock01_0 m3_12480_15420# m3_12480_15420# m1_15020_16390# m3_12560_15140# m1_14500_16280#
+ w_n610_16180# block01
Xnmos_08_0 m3_n5550_10400# cs_p_5_0/Vb cap_1/VSUBS cap_1/VSUBS nmos_08
Xblock0102_0 m1_14500_16280# m1_15020_16390# cap_1/VSUBS m1_20250_14460# block02
Xcap_1 m1_15020_16390# m3_12480_15420# m1_14500_16280# m3_12560_15140# cap_1/VSUBS
+ cap
Xres_0 m1_14500_16280# m1_15020_16390# m1_23690_16420# res
Xblock04_0 Diff_opamp_ly_0/diff_in_04_0/Vref m3_17920_18750# m1_20250_14460# m1_23690_16420#
+ m1_20250_14460# m1_20390_14580# w_n610_16180# block04
Xswitchblock_1 switchblock_1/beta bias_dummy_0/Vbias1 bias_dummy_0/Vbias2 bias_dummy_0/Vbias3
+ bias_dummy_0/Vbias4 switchblock_1/en_1 switchblock_1/en_2 m1_n7370_12690# m3_n7330_11130#
+ m1_n7650_12630# m3_n5550_10400# cap_1/VSUBS w_n610_16180# m1_n9150_12330# m1_n9750_12240#
+ m1_n8550_12540# Diff_opamp_ly_0/Vbias2 Diff_opamp_ly_0/Vbias3 Diff_opamp_ly_0/nmos_cload_01_1/Vbias1
+ switchblock
Xswitchblock_0 w_n610_16180# m1_n9750_12240# m1_n9150_12330# m1_n7650_12630# m1_n8550_12540#
+ m1_n7370_12690# switchblock01
Xbias_dummy_0 bias_dummy_0/Vbias1 bias_dummy_0/Vbias2 bias_dummy_0/Vbias3 bias_dummy_0/Vbias4
+ switchblock_1/beta cap_1/VSUBS cap_1/VSUBS bias_dummy_0/PBias w_n610_16180# bias_dummy
XDiff_opamp_ly_0 Diff_opamp_ly_0/Vbias3 Diff_opamp_ly_0/Vbias2 cap_1/VSUBS Diff_opamp_ly_0/nmos_cload_01_1/Vbias1
+ m3_12560_15140# cap_1/VSUBS Diff_opamp_ly_0/diff_in_04_0/Vref cap_1/VSUBS cap_1/VSUBS
+ cap_1/VSUBS cap_1/VSUBS cap_1/VSUBS Diff_opamp_ly_0/diff_in_03_0/in- cap_1/VSUBS
+ cap_1/VSUBS Diff_opamp_ly_0/li_12480_21783# Diff_opamp_ly_0/nmos_cload_01_1/a_n370_n2650#
+ m3_12480_15420# Diff_opamp_ly_0/diff_in_03_0/in+ cap_1/VSUBS Diff_opamp_ly_0/w_12480_21783#
+ m3_12480_15420# w_n610_16180# cap_1/VSUBS cap_1/VSUBS m3_n5550_10400# w_n610_16180#
+ Diff_opamp_ly
.ends

.subckt op_amp_lvs_final Rgm Vop Vm en_1 Vdd Vss Vref en_2 Vom Vp
X2stage_op_amp_1 Vop Vdd Rgm en_2 en_2 en_1 Vdd 2stage_op_amp_1/bias_dummy_0/PBias
+ Vom Vp Vdd Vdd Vref Vm Vdd Vss Vdd en_1 Vom Vdd Vss x2stage_op_amp
.ends

