magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect 5637 24985 10413 25073
rect 5637 13430 5673 24985
rect 5707 23223 10413 24985
rect 5707 23187 11283 23223
rect 23277 23187 34373 23223
rect 5707 23153 11373 23187
rect 23277 23180 23960 23187
rect 5707 21848 11283 23153
rect 5707 16567 10343 21848
rect 10377 16567 11283 21848
rect 23277 23137 23313 23180
rect 23347 23153 23960 23180
rect 33930 23153 34373 23187
rect 23347 23137 34373 23153
rect 23277 22700 34373 23137
rect 5707 16533 11342 16567
rect 5707 13430 10343 16533
rect 5637 13243 10343 13430
rect 10377 16497 11283 16533
rect 23277 16530 23313 22700
rect 23347 16530 34373 22700
rect 23277 16497 34373 16530
rect 10377 13243 10413 16497
rect 5637 13207 10413 13243
<< pwell >>
rect 547 20927 5223 21013
rect 547 11583 633 20927
rect 5137 11583 5223 20927
rect 34554 16374 34736 16556
rect 547 11497 5223 11583
<< psubdiff >>
rect 573 20953 658 20987
rect 692 20953 726 20987
rect 760 20953 794 20987
rect 828 20953 862 20987
rect 896 20953 930 20987
rect 964 20953 998 20987
rect 1032 20953 1066 20987
rect 1100 20953 1134 20987
rect 1168 20953 1202 20987
rect 1236 20953 1270 20987
rect 1304 20953 1338 20987
rect 1372 20953 1406 20987
rect 1440 20953 1474 20987
rect 1508 20953 1542 20987
rect 1576 20953 1610 20987
rect 1644 20953 1678 20987
rect 1712 20953 1746 20987
rect 1780 20953 1814 20987
rect 1848 20953 1882 20987
rect 1916 20953 1950 20987
rect 1984 20953 2018 20987
rect 2052 20953 2086 20987
rect 2120 20953 2154 20987
rect 2188 20953 2222 20987
rect 2256 20953 2290 20987
rect 2324 20953 2358 20987
rect 2392 20953 2426 20987
rect 2460 20953 2494 20987
rect 2528 20953 2562 20987
rect 2596 20953 2630 20987
rect 2664 20953 2698 20987
rect 2732 20953 2766 20987
rect 2800 20953 2834 20987
rect 2868 20953 2902 20987
rect 2936 20953 2970 20987
rect 3004 20953 3038 20987
rect 3072 20953 3106 20987
rect 3140 20953 3174 20987
rect 3208 20953 3242 20987
rect 3276 20953 3310 20987
rect 3344 20953 3378 20987
rect 3412 20953 3446 20987
rect 3480 20953 3514 20987
rect 3548 20953 3582 20987
rect 3616 20953 3650 20987
rect 3684 20953 3718 20987
rect 3752 20953 3786 20987
rect 3820 20953 3854 20987
rect 3888 20953 3922 20987
rect 3956 20953 3990 20987
rect 4024 20953 4058 20987
rect 4092 20953 4126 20987
rect 4160 20953 4194 20987
rect 4228 20953 4262 20987
rect 4296 20953 4330 20987
rect 4364 20953 4398 20987
rect 4432 20953 4466 20987
rect 4500 20953 4534 20987
rect 4568 20953 4602 20987
rect 4636 20953 4670 20987
rect 4704 20953 4738 20987
rect 4772 20953 4806 20987
rect 4840 20953 4874 20987
rect 4908 20953 4942 20987
rect 4976 20953 5010 20987
rect 5044 20953 5078 20987
rect 5112 20953 5197 20987
rect 573 20896 607 20953
rect 573 20828 607 20862
rect 573 20760 607 20794
rect 573 20692 607 20726
rect 573 20624 607 20658
rect 573 20556 607 20590
rect 573 20488 607 20522
rect 573 20420 607 20454
rect 573 20352 607 20386
rect 573 20284 607 20318
rect 573 20216 607 20250
rect 573 20148 607 20182
rect 573 20080 607 20114
rect 573 20012 607 20046
rect 573 19944 607 19978
rect 573 19876 607 19910
rect 573 19808 607 19842
rect 573 19740 607 19774
rect 573 19672 607 19706
rect 573 19604 607 19638
rect 573 19536 607 19570
rect 573 19468 607 19502
rect 573 19400 607 19434
rect 573 19332 607 19366
rect 573 19264 607 19298
rect 573 19196 607 19230
rect 573 19128 607 19162
rect 573 19060 607 19094
rect 573 18992 607 19026
rect 573 18924 607 18958
rect 573 18856 607 18890
rect 573 18788 607 18822
rect 573 18720 607 18754
rect 573 18652 607 18686
rect 573 18584 607 18618
rect 573 18516 607 18550
rect 573 18448 607 18482
rect 573 18380 607 18414
rect 573 18312 607 18346
rect 573 18244 607 18278
rect 573 18176 607 18210
rect 573 18108 607 18142
rect 573 18040 607 18074
rect 573 17972 607 18006
rect 573 17904 607 17938
rect 573 17836 607 17870
rect 573 17768 607 17802
rect 573 17700 607 17734
rect 573 17632 607 17666
rect 573 17564 607 17598
rect 573 17496 607 17530
rect 573 17428 607 17462
rect 573 17360 607 17394
rect 573 17292 607 17326
rect 573 17224 607 17258
rect 573 17156 607 17190
rect 573 17088 607 17122
rect 573 17020 607 17054
rect 573 16952 607 16986
rect 573 16884 607 16918
rect 573 16816 607 16850
rect 573 16748 607 16782
rect 573 16680 607 16714
rect 573 16612 607 16646
rect 573 16544 607 16578
rect 573 16476 607 16510
rect 573 16408 607 16442
rect 573 16340 607 16374
rect 573 16272 607 16306
rect 573 16204 607 16238
rect 573 16136 607 16170
rect 573 16068 607 16102
rect 573 16000 607 16034
rect 573 15932 607 15966
rect 573 15864 607 15898
rect 573 15796 607 15830
rect 573 15728 607 15762
rect 573 15660 607 15694
rect 573 15592 607 15626
rect 573 15524 607 15558
rect 573 15456 607 15490
rect 573 15388 607 15422
rect 573 15320 607 15354
rect 573 15252 607 15286
rect 573 15184 607 15218
rect 573 15116 607 15150
rect 573 15048 607 15082
rect 573 14980 607 15014
rect 573 14912 607 14946
rect 573 14844 607 14878
rect 573 14776 607 14810
rect 573 14708 607 14742
rect 573 14640 607 14674
rect 573 14572 607 14606
rect 573 14504 607 14538
rect 573 14436 607 14470
rect 573 14368 607 14402
rect 573 14300 607 14334
rect 573 14232 607 14266
rect 573 14164 607 14198
rect 573 14096 607 14130
rect 573 14028 607 14062
rect 573 13960 607 13994
rect 573 13892 607 13926
rect 573 13824 607 13858
rect 573 13756 607 13790
rect 573 13688 607 13722
rect 573 13620 607 13654
rect 573 13552 607 13586
rect 573 13484 607 13518
rect 573 13416 607 13450
rect 573 13348 607 13382
rect 573 13280 607 13314
rect 573 13212 607 13246
rect 573 13144 607 13178
rect 573 13076 607 13110
rect 573 13008 607 13042
rect 573 12940 607 12974
rect 573 12872 607 12906
rect 573 12804 607 12838
rect 573 12736 607 12770
rect 573 12668 607 12702
rect 573 12600 607 12634
rect 573 12532 607 12566
rect 573 12464 607 12498
rect 573 12396 607 12430
rect 573 12328 607 12362
rect 573 12260 607 12294
rect 573 12192 607 12226
rect 573 12124 607 12158
rect 573 12056 607 12090
rect 573 11988 607 12022
rect 573 11920 607 11954
rect 573 11852 607 11886
rect 573 11784 607 11818
rect 573 11716 607 11750
rect 573 11648 607 11682
rect 573 11557 607 11614
rect 5163 20896 5197 20953
rect 5163 20828 5197 20862
rect 5163 20760 5197 20794
rect 5163 20692 5197 20726
rect 5163 20624 5197 20658
rect 5163 20556 5197 20590
rect 5163 20488 5197 20522
rect 5163 20420 5197 20454
rect 5163 20352 5197 20386
rect 5163 20284 5197 20318
rect 5163 20216 5197 20250
rect 5163 20148 5197 20182
rect 5163 20080 5197 20114
rect 5163 20012 5197 20046
rect 5163 19944 5197 19978
rect 5163 19876 5197 19910
rect 5163 19808 5197 19842
rect 5163 19740 5197 19774
rect 5163 19672 5197 19706
rect 5163 19604 5197 19638
rect 5163 19536 5197 19570
rect 5163 19468 5197 19502
rect 5163 19400 5197 19434
rect 5163 19332 5197 19366
rect 5163 19264 5197 19298
rect 5163 19196 5197 19230
rect 5163 19128 5197 19162
rect 5163 19060 5197 19094
rect 5163 18992 5197 19026
rect 5163 18924 5197 18958
rect 5163 18856 5197 18890
rect 5163 18788 5197 18822
rect 5163 18720 5197 18754
rect 5163 18652 5197 18686
rect 5163 18584 5197 18618
rect 5163 18516 5197 18550
rect 5163 18448 5197 18482
rect 5163 18380 5197 18414
rect 5163 18312 5197 18346
rect 5163 18244 5197 18278
rect 5163 18176 5197 18210
rect 5163 18108 5197 18142
rect 5163 18040 5197 18074
rect 5163 17972 5197 18006
rect 5163 17904 5197 17938
rect 5163 17836 5197 17870
rect 5163 17768 5197 17802
rect 5163 17700 5197 17734
rect 5163 17632 5197 17666
rect 5163 17564 5197 17598
rect 5163 17496 5197 17530
rect 5163 17428 5197 17462
rect 5163 17360 5197 17394
rect 5163 17292 5197 17326
rect 5163 17224 5197 17258
rect 5163 17156 5197 17190
rect 5163 17088 5197 17122
rect 5163 17020 5197 17054
rect 5163 16952 5197 16986
rect 5163 16884 5197 16918
rect 5163 16816 5197 16850
rect 5163 16748 5197 16782
rect 5163 16680 5197 16714
rect 5163 16612 5197 16646
rect 5163 16544 5197 16578
rect 5163 16476 5197 16510
rect 5163 16408 5197 16442
rect 5163 16340 5197 16374
rect 5163 16272 5197 16306
rect 5163 16204 5197 16238
rect 5163 16136 5197 16170
rect 5163 16068 5197 16102
rect 5163 16000 5197 16034
rect 5163 15932 5197 15966
rect 5163 15864 5197 15898
rect 5163 15796 5197 15830
rect 5163 15728 5197 15762
rect 5163 15660 5197 15694
rect 5163 15592 5197 15626
rect 5163 15524 5197 15558
rect 5163 15456 5197 15490
rect 5163 15388 5197 15422
rect 5163 15320 5197 15354
rect 5163 15252 5197 15286
rect 5163 15184 5197 15218
rect 5163 15116 5197 15150
rect 5163 15048 5197 15082
rect 5163 14980 5197 15014
rect 5163 14912 5197 14946
rect 5163 14844 5197 14878
rect 5163 14776 5197 14810
rect 5163 14708 5197 14742
rect 5163 14640 5197 14674
rect 5163 14572 5197 14606
rect 5163 14504 5197 14538
rect 5163 14436 5197 14470
rect 5163 14368 5197 14402
rect 5163 14300 5197 14334
rect 5163 14232 5197 14266
rect 5163 14164 5197 14198
rect 5163 14096 5197 14130
rect 5163 14028 5197 14062
rect 5163 13960 5197 13994
rect 5163 13892 5197 13926
rect 5163 13824 5197 13858
rect 5163 13756 5197 13790
rect 5163 13688 5197 13722
rect 5163 13620 5197 13654
rect 5163 13552 5197 13586
rect 5163 13484 5197 13518
rect 5163 13416 5197 13450
rect 5163 13348 5197 13382
rect 5163 13280 5197 13314
rect 5163 13212 5197 13246
rect 34580 16447 34710 16530
rect 34580 16413 34623 16447
rect 34657 16413 34710 16447
rect 34580 16400 34710 16413
rect 5163 13144 5197 13178
rect 5163 13076 5197 13110
rect 5163 13008 5197 13042
rect 5163 12940 5197 12974
rect 5163 12872 5197 12906
rect 5163 12804 5197 12838
rect 5163 12736 5197 12770
rect 5163 12668 5197 12702
rect 5163 12600 5197 12634
rect 5163 12532 5197 12566
rect 5163 12464 5197 12498
rect 5163 12396 5197 12430
rect 5163 12328 5197 12362
rect 5163 12260 5197 12294
rect 5163 12192 5197 12226
rect 5163 12124 5197 12158
rect 5163 12056 5197 12090
rect 5163 11988 5197 12022
rect 5163 11920 5197 11954
rect 5163 11852 5197 11886
rect 5163 11784 5197 11818
rect 5163 11716 5197 11750
rect 5163 11648 5197 11682
rect 5163 11557 5197 11614
rect 573 11523 658 11557
rect 692 11523 726 11557
rect 760 11523 794 11557
rect 828 11523 862 11557
rect 896 11523 930 11557
rect 964 11523 998 11557
rect 1032 11523 1066 11557
rect 1100 11523 1134 11557
rect 1168 11523 1202 11557
rect 1236 11523 1270 11557
rect 1304 11523 1338 11557
rect 1372 11523 1406 11557
rect 1440 11523 1474 11557
rect 1508 11523 1542 11557
rect 1576 11523 1610 11557
rect 1644 11523 1678 11557
rect 1712 11523 1746 11557
rect 1780 11523 1814 11557
rect 1848 11523 1882 11557
rect 1916 11523 1950 11557
rect 1984 11523 2018 11557
rect 2052 11523 2086 11557
rect 2120 11523 2154 11557
rect 2188 11523 2222 11557
rect 2256 11523 2290 11557
rect 2324 11523 2358 11557
rect 2392 11523 2426 11557
rect 2460 11523 2494 11557
rect 2528 11523 2562 11557
rect 2596 11523 2630 11557
rect 2664 11523 2698 11557
rect 2732 11523 2766 11557
rect 2800 11523 2834 11557
rect 2868 11523 2902 11557
rect 2936 11523 2970 11557
rect 3004 11523 3038 11557
rect 3072 11523 3106 11557
rect 3140 11523 3174 11557
rect 3208 11523 3242 11557
rect 3276 11523 3310 11557
rect 3344 11523 3378 11557
rect 3412 11523 3446 11557
rect 3480 11523 3514 11557
rect 3548 11523 3582 11557
rect 3616 11523 3650 11557
rect 3684 11523 3718 11557
rect 3752 11523 3786 11557
rect 3820 11523 3854 11557
rect 3888 11523 3922 11557
rect 3956 11523 3990 11557
rect 4024 11523 4058 11557
rect 4092 11523 4126 11557
rect 4160 11523 4194 11557
rect 4228 11523 4262 11557
rect 4296 11523 4330 11557
rect 4364 11523 4398 11557
rect 4432 11523 4466 11557
rect 4500 11523 4534 11557
rect 4568 11523 4602 11557
rect 4636 11523 4670 11557
rect 4704 11523 4738 11557
rect 4772 11523 4806 11557
rect 4840 11523 4874 11557
rect 4908 11523 4942 11557
rect 4976 11523 5010 11557
rect 5044 11523 5078 11557
rect 5112 11523 5197 11557
<< nsubdiff >>
rect 5673 25003 5764 25037
rect 5798 25003 5832 25037
rect 5866 25003 5900 25037
rect 5934 25003 5968 25037
rect 6002 25003 6036 25037
rect 6070 25003 6104 25037
rect 6138 25003 6172 25037
rect 6206 25003 6240 25037
rect 6274 25003 6308 25037
rect 6342 25003 6376 25037
rect 6410 25003 6444 25037
rect 6478 25003 6512 25037
rect 6546 25003 6580 25037
rect 6614 25003 6648 25037
rect 6682 25003 6716 25037
rect 6750 25003 6784 25037
rect 6818 25003 6852 25037
rect 6886 25003 6920 25037
rect 6954 25003 6988 25037
rect 7022 25003 7056 25037
rect 7090 25003 7124 25037
rect 7158 25003 7192 25037
rect 7226 25003 7260 25037
rect 7294 25003 7328 25037
rect 7362 25003 7396 25037
rect 7430 25003 7464 25037
rect 7498 25003 7532 25037
rect 7566 25003 7600 25037
rect 7634 25003 7668 25037
rect 7702 25003 7736 25037
rect 7770 25003 7804 25037
rect 7838 25003 7872 25037
rect 7906 25003 7940 25037
rect 7974 25003 8008 25037
rect 8042 25003 8076 25037
rect 8110 25003 8144 25037
rect 8178 25003 8212 25037
rect 8246 25003 8280 25037
rect 8314 25003 8348 25037
rect 8382 25003 8416 25037
rect 8450 25003 8484 25037
rect 8518 25003 8552 25037
rect 8586 25003 8620 25037
rect 8654 25003 8688 25037
rect 8722 25003 8756 25037
rect 8790 25003 8824 25037
rect 8858 25003 8892 25037
rect 8926 25003 8960 25037
rect 8994 25003 9028 25037
rect 9062 25003 9096 25037
rect 9130 25003 9164 25037
rect 9198 25003 9232 25037
rect 9266 25003 9300 25037
rect 9334 25003 9368 25037
rect 9402 25003 9436 25037
rect 9470 25003 9504 25037
rect 9538 25003 9572 25037
rect 9606 25003 9640 25037
rect 9674 25003 9708 25037
rect 9742 25003 9776 25037
rect 9810 25003 9844 25037
rect 9878 25003 9912 25037
rect 9946 25003 9980 25037
rect 10014 25003 10048 25037
rect 10082 25003 10116 25037
rect 10150 25003 10184 25037
rect 10218 25003 10252 25037
rect 10286 25003 10377 25037
rect 5673 24985 5707 25003
rect 10343 24947 10377 25003
rect 10343 24879 10377 24913
rect 10343 24811 10377 24845
rect 10343 24743 10377 24777
rect 10343 24675 10377 24709
rect 10343 24607 10377 24641
rect 10343 24539 10377 24573
rect 10343 24471 10377 24505
rect 10343 24403 10377 24437
rect 10343 24335 10377 24369
rect 10343 24267 10377 24301
rect 10343 24199 10377 24233
rect 10343 24131 10377 24165
rect 10343 24063 10377 24097
rect 10343 23995 10377 24029
rect 10343 23927 10377 23961
rect 10343 23859 10377 23893
rect 10343 23187 10377 23825
rect 10343 23153 11373 23187
rect 23313 23180 23426 23187
rect 23347 23153 23426 23180
rect 23460 23153 23494 23187
rect 23528 23153 23562 23187
rect 23596 23153 23630 23187
rect 23664 23153 23698 23187
rect 23732 23153 23766 23187
rect 23800 23153 23960 23187
rect 33930 23153 34078 23187
rect 34112 23153 34146 23187
rect 34180 23153 34214 23187
rect 34248 23153 34337 23187
rect 10343 21882 10377 23153
rect 23313 22700 23347 23137
rect 34303 23107 34337 23153
rect 34303 23039 34337 23073
rect 34303 22971 34337 23005
rect 34303 22903 34337 22937
rect 34303 22835 34337 22869
rect 34303 22767 34337 22801
rect 10308 21848 10377 21882
rect 34303 22699 34337 22733
rect 34303 22631 34337 22665
rect 34303 22563 34337 22597
rect 34303 22495 34337 22529
rect 34303 22427 34337 22461
rect 34303 22359 34337 22393
rect 34303 22291 34337 22325
rect 34303 22223 34337 22257
rect 34303 22155 34337 22189
rect 34303 22087 34337 22121
rect 34303 22019 34337 22053
rect 34303 21951 34337 21985
rect 34303 21883 34337 21917
rect 34303 21815 34337 21849
rect 34303 21747 34337 21781
rect 34303 21679 34337 21713
rect 34303 21611 34337 21645
rect 34303 21543 34337 21577
rect 34303 21475 34337 21509
rect 34303 21407 34337 21441
rect 34303 21339 34337 21373
rect 34303 21271 34337 21305
rect 34303 21203 34337 21237
rect 34303 21135 34337 21169
rect 34303 21067 34337 21101
rect 34303 20999 34337 21033
rect 34303 20931 34337 20965
rect 34303 20863 34337 20897
rect 34303 20795 34337 20829
rect 34303 20727 34337 20761
rect 34303 20659 34337 20693
rect 34303 20591 34337 20625
rect 34303 20523 34337 20557
rect 34303 20455 34337 20489
rect 34303 20387 34337 20421
rect 34303 20319 34337 20353
rect 34303 20251 34337 20285
rect 34303 20183 34337 20217
rect 34303 20115 34337 20149
rect 34303 20047 34337 20081
rect 34303 19979 34337 20013
rect 34303 19911 34337 19945
rect 34303 19843 34337 19877
rect 34303 19775 34337 19809
rect 34303 19707 34337 19741
rect 34303 19639 34337 19673
rect 34303 19571 34337 19605
rect 34303 19503 34337 19537
rect 34303 19435 34337 19469
rect 34303 19367 34337 19401
rect 34303 19299 34337 19333
rect 34303 19231 34337 19265
rect 34303 19163 34337 19197
rect 34303 19095 34337 19129
rect 34303 19027 34337 19061
rect 34303 18959 34337 18993
rect 34303 18891 34337 18925
rect 34303 18823 34337 18857
rect 34303 18755 34337 18789
rect 34303 18687 34337 18721
rect 34303 18619 34337 18653
rect 34303 18551 34337 18585
rect 10320 16567 10343 18523
rect 34303 18483 34337 18517
rect 34303 18415 34337 18449
rect 34303 18347 34337 18381
rect 34303 18279 34337 18313
rect 34303 18211 34337 18245
rect 34303 18143 34337 18177
rect 34303 18075 34337 18109
rect 34303 18007 34337 18041
rect 34303 17939 34337 17973
rect 34303 17871 34337 17905
rect 34303 17803 34337 17837
rect 34303 17735 34337 17769
rect 34303 17667 34337 17701
rect 34303 17599 34337 17633
rect 34303 17531 34337 17565
rect 34303 17463 34337 17497
rect 34303 17395 34337 17429
rect 34303 17327 34337 17361
rect 34303 17259 34337 17293
rect 34303 17191 34337 17225
rect 34303 17123 34337 17157
rect 34303 17055 34337 17089
rect 34303 16987 34337 17021
rect 34303 16919 34337 16953
rect 34303 16851 34337 16885
rect 34303 16783 34337 16817
rect 34303 16715 34337 16749
rect 34303 16647 34337 16681
rect 34303 16567 34337 16613
rect 10320 16533 11342 16567
rect 23347 16533 23417 16567
rect 23451 16533 23485 16567
rect 23519 16533 23553 16567
rect 23587 16533 23621 16567
rect 23655 16533 23689 16567
rect 23723 16533 23757 16567
rect 23791 16533 23825 16567
rect 23859 16533 23893 16567
rect 23927 16533 23961 16567
rect 23995 16533 24029 16567
rect 24063 16533 24097 16567
rect 24131 16533 24165 16567
rect 24199 16533 24233 16567
rect 24267 16533 24301 16567
rect 24335 16533 24369 16567
rect 24403 16533 24437 16567
rect 24471 16533 24505 16567
rect 24539 16533 24573 16567
rect 24607 16533 24641 16567
rect 24675 16533 24709 16567
rect 24743 16533 24777 16567
rect 24811 16533 24845 16567
rect 24879 16533 24913 16567
rect 24947 16533 24981 16567
rect 25015 16533 25049 16567
rect 25083 16533 25117 16567
rect 25151 16533 25185 16567
rect 25219 16533 25253 16567
rect 25287 16533 25321 16567
rect 25355 16533 25389 16567
rect 25423 16533 25457 16567
rect 25491 16533 25525 16567
rect 25559 16533 25593 16567
rect 25627 16533 25661 16567
rect 25695 16533 25729 16567
rect 25763 16533 25797 16567
rect 25831 16533 25865 16567
rect 25899 16533 25933 16567
rect 25967 16533 26001 16567
rect 26035 16533 26069 16567
rect 26103 16533 26137 16567
rect 26171 16533 26205 16567
rect 26239 16533 26273 16567
rect 26307 16533 26341 16567
rect 26375 16533 26409 16567
rect 26443 16533 26477 16567
rect 26511 16533 26545 16567
rect 26579 16533 26613 16567
rect 26647 16533 26681 16567
rect 26715 16533 26749 16567
rect 26783 16533 26817 16567
rect 26851 16533 26885 16567
rect 26919 16533 26953 16567
rect 26987 16533 27021 16567
rect 27055 16533 27089 16567
rect 27123 16533 27157 16567
rect 27191 16533 27225 16567
rect 27259 16533 27293 16567
rect 27327 16533 27361 16567
rect 27395 16533 27429 16567
rect 27463 16533 27497 16567
rect 27531 16533 27565 16567
rect 27599 16533 27633 16567
rect 27667 16533 27701 16567
rect 27735 16533 27769 16567
rect 27803 16533 27837 16567
rect 27871 16533 27905 16567
rect 27939 16533 27973 16567
rect 28007 16533 28041 16567
rect 28075 16533 28109 16567
rect 28143 16533 28177 16567
rect 28211 16533 28245 16567
rect 28279 16533 28313 16567
rect 28347 16533 28381 16567
rect 28415 16533 28449 16567
rect 28483 16533 28517 16567
rect 28551 16533 28585 16567
rect 28619 16533 28653 16567
rect 28687 16533 28721 16567
rect 28755 16533 28789 16567
rect 28823 16533 28857 16567
rect 28891 16533 28925 16567
rect 28959 16533 28993 16567
rect 29027 16533 29061 16567
rect 29095 16533 29129 16567
rect 29163 16533 29197 16567
rect 29231 16533 29265 16567
rect 29299 16533 29333 16567
rect 29367 16533 29401 16567
rect 29435 16533 29469 16567
rect 29503 16533 29537 16567
rect 29571 16533 29605 16567
rect 29639 16533 29673 16567
rect 29707 16533 29741 16567
rect 29775 16533 29809 16567
rect 29843 16533 29877 16567
rect 29911 16533 29945 16567
rect 29979 16533 30013 16567
rect 30047 16533 30081 16567
rect 30115 16533 30149 16567
rect 30183 16533 30217 16567
rect 30251 16533 30285 16567
rect 30319 16533 30353 16567
rect 30387 16533 30421 16567
rect 30455 16533 30489 16567
rect 30523 16533 30557 16567
rect 30591 16533 30625 16567
rect 30659 16533 30693 16567
rect 30727 16533 30761 16567
rect 30795 16533 30829 16567
rect 30863 16533 30897 16567
rect 30931 16533 30965 16567
rect 30999 16533 31033 16567
rect 31067 16533 31101 16567
rect 31135 16533 31169 16567
rect 31203 16533 31237 16567
rect 31271 16533 31305 16567
rect 31339 16533 31373 16567
rect 31407 16533 31441 16567
rect 31475 16533 31509 16567
rect 31543 16533 31577 16567
rect 31611 16533 31645 16567
rect 31679 16533 31713 16567
rect 31747 16533 31781 16567
rect 31815 16533 31849 16567
rect 31883 16533 31917 16567
rect 31951 16533 31985 16567
rect 32019 16533 32053 16567
rect 32087 16533 32121 16567
rect 32155 16533 32189 16567
rect 32223 16533 32257 16567
rect 32291 16533 32325 16567
rect 32359 16533 32393 16567
rect 32427 16533 32461 16567
rect 32495 16533 32529 16567
rect 32563 16533 32597 16567
rect 32631 16533 32665 16567
rect 32699 16533 32733 16567
rect 32767 16533 32801 16567
rect 32835 16533 32869 16567
rect 32903 16533 32937 16567
rect 32971 16533 33005 16567
rect 33039 16533 33073 16567
rect 33107 16533 33141 16567
rect 33175 16533 33209 16567
rect 33243 16533 33277 16567
rect 33311 16533 33345 16567
rect 33379 16533 33413 16567
rect 33447 16533 33481 16567
rect 33515 16533 33549 16567
rect 33583 16533 33617 16567
rect 33651 16533 33685 16567
rect 33719 16533 33753 16567
rect 33787 16533 33821 16567
rect 33855 16533 33889 16567
rect 33923 16533 33957 16567
rect 33991 16533 34025 16567
rect 34059 16533 34093 16567
rect 34127 16533 34161 16567
rect 34195 16533 34229 16567
rect 34263 16533 34337 16567
rect 5673 13396 5744 13430
rect 5673 13367 5707 13396
rect 5673 13277 5707 13333
rect 10320 13330 10343 16533
rect 10310 13277 10343 13330
rect 5673 13243 5764 13277
rect 5798 13243 5832 13277
rect 5866 13243 5900 13277
rect 5934 13243 5968 13277
rect 6002 13243 6036 13277
rect 6070 13243 6104 13277
rect 6138 13243 6172 13277
rect 6206 13243 6240 13277
rect 6274 13243 6308 13277
rect 6342 13243 6376 13277
rect 6410 13243 6444 13277
rect 6478 13243 6512 13277
rect 6546 13243 6580 13277
rect 6614 13243 6648 13277
rect 6682 13243 6716 13277
rect 6750 13243 6784 13277
rect 6818 13243 6852 13277
rect 6886 13243 6920 13277
rect 6954 13243 6988 13277
rect 7022 13243 7056 13277
rect 7090 13243 7124 13277
rect 7158 13243 7192 13277
rect 7226 13243 7260 13277
rect 7294 13243 7328 13277
rect 7362 13243 7396 13277
rect 7430 13243 7464 13277
rect 7498 13243 7532 13277
rect 7566 13243 7600 13277
rect 7634 13243 7668 13277
rect 7702 13243 7736 13277
rect 7770 13243 7804 13277
rect 7838 13243 7872 13277
rect 7906 13243 7940 13277
rect 7974 13243 8008 13277
rect 8042 13243 8076 13277
rect 8110 13243 8144 13277
rect 8178 13243 8212 13277
rect 8246 13243 8280 13277
rect 8314 13243 8348 13277
rect 8382 13243 8416 13277
rect 8450 13243 8484 13277
rect 8518 13243 8552 13277
rect 8586 13243 8620 13277
rect 8654 13243 8688 13277
rect 8722 13243 8756 13277
rect 8790 13243 8824 13277
rect 8858 13243 8892 13277
rect 8926 13243 8960 13277
rect 8994 13243 9028 13277
rect 9062 13243 9096 13277
rect 9130 13243 9164 13277
rect 9198 13243 9232 13277
rect 9266 13243 9300 13277
rect 9334 13243 9368 13277
rect 9402 13243 9436 13277
rect 9470 13243 9504 13277
rect 9538 13243 9572 13277
rect 9606 13243 9640 13277
rect 9674 13243 9708 13277
rect 9742 13243 9776 13277
rect 9810 13243 9844 13277
rect 9878 13243 9912 13277
rect 9946 13243 9980 13277
rect 10014 13243 10048 13277
rect 10082 13243 10116 13277
rect 10150 13243 10184 13277
rect 10218 13243 10252 13277
rect 10286 13243 10343 13277
<< psubdiffcont >>
rect 658 20953 692 20987
rect 726 20953 760 20987
rect 794 20953 828 20987
rect 862 20953 896 20987
rect 930 20953 964 20987
rect 998 20953 1032 20987
rect 1066 20953 1100 20987
rect 1134 20953 1168 20987
rect 1202 20953 1236 20987
rect 1270 20953 1304 20987
rect 1338 20953 1372 20987
rect 1406 20953 1440 20987
rect 1474 20953 1508 20987
rect 1542 20953 1576 20987
rect 1610 20953 1644 20987
rect 1678 20953 1712 20987
rect 1746 20953 1780 20987
rect 1814 20953 1848 20987
rect 1882 20953 1916 20987
rect 1950 20953 1984 20987
rect 2018 20953 2052 20987
rect 2086 20953 2120 20987
rect 2154 20953 2188 20987
rect 2222 20953 2256 20987
rect 2290 20953 2324 20987
rect 2358 20953 2392 20987
rect 2426 20953 2460 20987
rect 2494 20953 2528 20987
rect 2562 20953 2596 20987
rect 2630 20953 2664 20987
rect 2698 20953 2732 20987
rect 2766 20953 2800 20987
rect 2834 20953 2868 20987
rect 2902 20953 2936 20987
rect 2970 20953 3004 20987
rect 3038 20953 3072 20987
rect 3106 20953 3140 20987
rect 3174 20953 3208 20987
rect 3242 20953 3276 20987
rect 3310 20953 3344 20987
rect 3378 20953 3412 20987
rect 3446 20953 3480 20987
rect 3514 20953 3548 20987
rect 3582 20953 3616 20987
rect 3650 20953 3684 20987
rect 3718 20953 3752 20987
rect 3786 20953 3820 20987
rect 3854 20953 3888 20987
rect 3922 20953 3956 20987
rect 3990 20953 4024 20987
rect 4058 20953 4092 20987
rect 4126 20953 4160 20987
rect 4194 20953 4228 20987
rect 4262 20953 4296 20987
rect 4330 20953 4364 20987
rect 4398 20953 4432 20987
rect 4466 20953 4500 20987
rect 4534 20953 4568 20987
rect 4602 20953 4636 20987
rect 4670 20953 4704 20987
rect 4738 20953 4772 20987
rect 4806 20953 4840 20987
rect 4874 20953 4908 20987
rect 4942 20953 4976 20987
rect 5010 20953 5044 20987
rect 5078 20953 5112 20987
rect 573 20862 607 20896
rect 573 20794 607 20828
rect 573 20726 607 20760
rect 573 20658 607 20692
rect 573 20590 607 20624
rect 573 20522 607 20556
rect 573 20454 607 20488
rect 573 20386 607 20420
rect 573 20318 607 20352
rect 573 20250 607 20284
rect 573 20182 607 20216
rect 573 20114 607 20148
rect 573 20046 607 20080
rect 573 19978 607 20012
rect 573 19910 607 19944
rect 573 19842 607 19876
rect 573 19774 607 19808
rect 573 19706 607 19740
rect 573 19638 607 19672
rect 573 19570 607 19604
rect 573 19502 607 19536
rect 573 19434 607 19468
rect 573 19366 607 19400
rect 573 19298 607 19332
rect 573 19230 607 19264
rect 573 19162 607 19196
rect 573 19094 607 19128
rect 573 19026 607 19060
rect 573 18958 607 18992
rect 573 18890 607 18924
rect 573 18822 607 18856
rect 573 18754 607 18788
rect 573 18686 607 18720
rect 573 18618 607 18652
rect 573 18550 607 18584
rect 573 18482 607 18516
rect 573 18414 607 18448
rect 573 18346 607 18380
rect 573 18278 607 18312
rect 573 18210 607 18244
rect 573 18142 607 18176
rect 573 18074 607 18108
rect 573 18006 607 18040
rect 573 17938 607 17972
rect 573 17870 607 17904
rect 573 17802 607 17836
rect 573 17734 607 17768
rect 573 17666 607 17700
rect 573 17598 607 17632
rect 573 17530 607 17564
rect 573 17462 607 17496
rect 573 17394 607 17428
rect 573 17326 607 17360
rect 573 17258 607 17292
rect 573 17190 607 17224
rect 573 17122 607 17156
rect 573 17054 607 17088
rect 573 16986 607 17020
rect 573 16918 607 16952
rect 573 16850 607 16884
rect 573 16782 607 16816
rect 573 16714 607 16748
rect 573 16646 607 16680
rect 573 16578 607 16612
rect 573 16510 607 16544
rect 573 16442 607 16476
rect 573 16374 607 16408
rect 573 16306 607 16340
rect 573 16238 607 16272
rect 573 16170 607 16204
rect 573 16102 607 16136
rect 573 16034 607 16068
rect 573 15966 607 16000
rect 573 15898 607 15932
rect 573 15830 607 15864
rect 573 15762 607 15796
rect 573 15694 607 15728
rect 573 15626 607 15660
rect 573 15558 607 15592
rect 573 15490 607 15524
rect 573 15422 607 15456
rect 573 15354 607 15388
rect 573 15286 607 15320
rect 573 15218 607 15252
rect 573 15150 607 15184
rect 573 15082 607 15116
rect 573 15014 607 15048
rect 573 14946 607 14980
rect 573 14878 607 14912
rect 573 14810 607 14844
rect 573 14742 607 14776
rect 573 14674 607 14708
rect 573 14606 607 14640
rect 573 14538 607 14572
rect 573 14470 607 14504
rect 573 14402 607 14436
rect 573 14334 607 14368
rect 573 14266 607 14300
rect 573 14198 607 14232
rect 573 14130 607 14164
rect 573 14062 607 14096
rect 573 13994 607 14028
rect 573 13926 607 13960
rect 573 13858 607 13892
rect 573 13790 607 13824
rect 573 13722 607 13756
rect 573 13654 607 13688
rect 573 13586 607 13620
rect 573 13518 607 13552
rect 573 13450 607 13484
rect 573 13382 607 13416
rect 573 13314 607 13348
rect 573 13246 607 13280
rect 573 13178 607 13212
rect 573 13110 607 13144
rect 573 13042 607 13076
rect 573 12974 607 13008
rect 573 12906 607 12940
rect 573 12838 607 12872
rect 573 12770 607 12804
rect 573 12702 607 12736
rect 573 12634 607 12668
rect 573 12566 607 12600
rect 573 12498 607 12532
rect 573 12430 607 12464
rect 573 12362 607 12396
rect 573 12294 607 12328
rect 573 12226 607 12260
rect 573 12158 607 12192
rect 573 12090 607 12124
rect 573 12022 607 12056
rect 573 11954 607 11988
rect 573 11886 607 11920
rect 573 11818 607 11852
rect 573 11750 607 11784
rect 573 11682 607 11716
rect 573 11614 607 11648
rect 5163 20862 5197 20896
rect 5163 20794 5197 20828
rect 5163 20726 5197 20760
rect 5163 20658 5197 20692
rect 5163 20590 5197 20624
rect 5163 20522 5197 20556
rect 5163 20454 5197 20488
rect 5163 20386 5197 20420
rect 5163 20318 5197 20352
rect 5163 20250 5197 20284
rect 5163 20182 5197 20216
rect 5163 20114 5197 20148
rect 5163 20046 5197 20080
rect 5163 19978 5197 20012
rect 5163 19910 5197 19944
rect 5163 19842 5197 19876
rect 5163 19774 5197 19808
rect 5163 19706 5197 19740
rect 5163 19638 5197 19672
rect 5163 19570 5197 19604
rect 5163 19502 5197 19536
rect 5163 19434 5197 19468
rect 5163 19366 5197 19400
rect 5163 19298 5197 19332
rect 5163 19230 5197 19264
rect 5163 19162 5197 19196
rect 5163 19094 5197 19128
rect 5163 19026 5197 19060
rect 5163 18958 5197 18992
rect 5163 18890 5197 18924
rect 5163 18822 5197 18856
rect 5163 18754 5197 18788
rect 5163 18686 5197 18720
rect 5163 18618 5197 18652
rect 5163 18550 5197 18584
rect 5163 18482 5197 18516
rect 5163 18414 5197 18448
rect 5163 18346 5197 18380
rect 5163 18278 5197 18312
rect 5163 18210 5197 18244
rect 5163 18142 5197 18176
rect 5163 18074 5197 18108
rect 5163 18006 5197 18040
rect 5163 17938 5197 17972
rect 5163 17870 5197 17904
rect 5163 17802 5197 17836
rect 5163 17734 5197 17768
rect 5163 17666 5197 17700
rect 5163 17598 5197 17632
rect 5163 17530 5197 17564
rect 5163 17462 5197 17496
rect 5163 17394 5197 17428
rect 5163 17326 5197 17360
rect 5163 17258 5197 17292
rect 5163 17190 5197 17224
rect 5163 17122 5197 17156
rect 5163 17054 5197 17088
rect 5163 16986 5197 17020
rect 5163 16918 5197 16952
rect 5163 16850 5197 16884
rect 5163 16782 5197 16816
rect 5163 16714 5197 16748
rect 5163 16646 5197 16680
rect 5163 16578 5197 16612
rect 5163 16510 5197 16544
rect 5163 16442 5197 16476
rect 5163 16374 5197 16408
rect 5163 16306 5197 16340
rect 5163 16238 5197 16272
rect 5163 16170 5197 16204
rect 5163 16102 5197 16136
rect 5163 16034 5197 16068
rect 5163 15966 5197 16000
rect 5163 15898 5197 15932
rect 5163 15830 5197 15864
rect 5163 15762 5197 15796
rect 5163 15694 5197 15728
rect 5163 15626 5197 15660
rect 5163 15558 5197 15592
rect 5163 15490 5197 15524
rect 5163 15422 5197 15456
rect 5163 15354 5197 15388
rect 5163 15286 5197 15320
rect 5163 15218 5197 15252
rect 5163 15150 5197 15184
rect 5163 15082 5197 15116
rect 5163 15014 5197 15048
rect 5163 14946 5197 14980
rect 5163 14878 5197 14912
rect 5163 14810 5197 14844
rect 5163 14742 5197 14776
rect 5163 14674 5197 14708
rect 5163 14606 5197 14640
rect 5163 14538 5197 14572
rect 5163 14470 5197 14504
rect 5163 14402 5197 14436
rect 5163 14334 5197 14368
rect 5163 14266 5197 14300
rect 5163 14198 5197 14232
rect 5163 14130 5197 14164
rect 5163 14062 5197 14096
rect 5163 13994 5197 14028
rect 5163 13926 5197 13960
rect 5163 13858 5197 13892
rect 5163 13790 5197 13824
rect 5163 13722 5197 13756
rect 5163 13654 5197 13688
rect 5163 13586 5197 13620
rect 5163 13518 5197 13552
rect 5163 13450 5197 13484
rect 5163 13382 5197 13416
rect 5163 13314 5197 13348
rect 5163 13246 5197 13280
rect 34623 16413 34657 16447
rect 5163 13178 5197 13212
rect 5163 13110 5197 13144
rect 5163 13042 5197 13076
rect 5163 12974 5197 13008
rect 5163 12906 5197 12940
rect 5163 12838 5197 12872
rect 5163 12770 5197 12804
rect 5163 12702 5197 12736
rect 5163 12634 5197 12668
rect 5163 12566 5197 12600
rect 5163 12498 5197 12532
rect 5163 12430 5197 12464
rect 5163 12362 5197 12396
rect 5163 12294 5197 12328
rect 5163 12226 5197 12260
rect 5163 12158 5197 12192
rect 5163 12090 5197 12124
rect 5163 12022 5197 12056
rect 5163 11954 5197 11988
rect 5163 11886 5197 11920
rect 5163 11818 5197 11852
rect 5163 11750 5197 11784
rect 5163 11682 5197 11716
rect 5163 11614 5197 11648
rect 658 11523 692 11557
rect 726 11523 760 11557
rect 794 11523 828 11557
rect 862 11523 896 11557
rect 930 11523 964 11557
rect 998 11523 1032 11557
rect 1066 11523 1100 11557
rect 1134 11523 1168 11557
rect 1202 11523 1236 11557
rect 1270 11523 1304 11557
rect 1338 11523 1372 11557
rect 1406 11523 1440 11557
rect 1474 11523 1508 11557
rect 1542 11523 1576 11557
rect 1610 11523 1644 11557
rect 1678 11523 1712 11557
rect 1746 11523 1780 11557
rect 1814 11523 1848 11557
rect 1882 11523 1916 11557
rect 1950 11523 1984 11557
rect 2018 11523 2052 11557
rect 2086 11523 2120 11557
rect 2154 11523 2188 11557
rect 2222 11523 2256 11557
rect 2290 11523 2324 11557
rect 2358 11523 2392 11557
rect 2426 11523 2460 11557
rect 2494 11523 2528 11557
rect 2562 11523 2596 11557
rect 2630 11523 2664 11557
rect 2698 11523 2732 11557
rect 2766 11523 2800 11557
rect 2834 11523 2868 11557
rect 2902 11523 2936 11557
rect 2970 11523 3004 11557
rect 3038 11523 3072 11557
rect 3106 11523 3140 11557
rect 3174 11523 3208 11557
rect 3242 11523 3276 11557
rect 3310 11523 3344 11557
rect 3378 11523 3412 11557
rect 3446 11523 3480 11557
rect 3514 11523 3548 11557
rect 3582 11523 3616 11557
rect 3650 11523 3684 11557
rect 3718 11523 3752 11557
rect 3786 11523 3820 11557
rect 3854 11523 3888 11557
rect 3922 11523 3956 11557
rect 3990 11523 4024 11557
rect 4058 11523 4092 11557
rect 4126 11523 4160 11557
rect 4194 11523 4228 11557
rect 4262 11523 4296 11557
rect 4330 11523 4364 11557
rect 4398 11523 4432 11557
rect 4466 11523 4500 11557
rect 4534 11523 4568 11557
rect 4602 11523 4636 11557
rect 4670 11523 4704 11557
rect 4738 11523 4772 11557
rect 4806 11523 4840 11557
rect 4874 11523 4908 11557
rect 4942 11523 4976 11557
rect 5010 11523 5044 11557
rect 5078 11523 5112 11557
<< nsubdiffcont >>
rect 5764 25003 5798 25037
rect 5832 25003 5866 25037
rect 5900 25003 5934 25037
rect 5968 25003 6002 25037
rect 6036 25003 6070 25037
rect 6104 25003 6138 25037
rect 6172 25003 6206 25037
rect 6240 25003 6274 25037
rect 6308 25003 6342 25037
rect 6376 25003 6410 25037
rect 6444 25003 6478 25037
rect 6512 25003 6546 25037
rect 6580 25003 6614 25037
rect 6648 25003 6682 25037
rect 6716 25003 6750 25037
rect 6784 25003 6818 25037
rect 6852 25003 6886 25037
rect 6920 25003 6954 25037
rect 6988 25003 7022 25037
rect 7056 25003 7090 25037
rect 7124 25003 7158 25037
rect 7192 25003 7226 25037
rect 7260 25003 7294 25037
rect 7328 25003 7362 25037
rect 7396 25003 7430 25037
rect 7464 25003 7498 25037
rect 7532 25003 7566 25037
rect 7600 25003 7634 25037
rect 7668 25003 7702 25037
rect 7736 25003 7770 25037
rect 7804 25003 7838 25037
rect 7872 25003 7906 25037
rect 7940 25003 7974 25037
rect 8008 25003 8042 25037
rect 8076 25003 8110 25037
rect 8144 25003 8178 25037
rect 8212 25003 8246 25037
rect 8280 25003 8314 25037
rect 8348 25003 8382 25037
rect 8416 25003 8450 25037
rect 8484 25003 8518 25037
rect 8552 25003 8586 25037
rect 8620 25003 8654 25037
rect 8688 25003 8722 25037
rect 8756 25003 8790 25037
rect 8824 25003 8858 25037
rect 8892 25003 8926 25037
rect 8960 25003 8994 25037
rect 9028 25003 9062 25037
rect 9096 25003 9130 25037
rect 9164 25003 9198 25037
rect 9232 25003 9266 25037
rect 9300 25003 9334 25037
rect 9368 25003 9402 25037
rect 9436 25003 9470 25037
rect 9504 25003 9538 25037
rect 9572 25003 9606 25037
rect 9640 25003 9674 25037
rect 9708 25003 9742 25037
rect 9776 25003 9810 25037
rect 9844 25003 9878 25037
rect 9912 25003 9946 25037
rect 9980 25003 10014 25037
rect 10048 25003 10082 25037
rect 10116 25003 10150 25037
rect 10184 25003 10218 25037
rect 10252 25003 10286 25037
rect 10343 24913 10377 24947
rect 10343 24845 10377 24879
rect 10343 24777 10377 24811
rect 10343 24709 10377 24743
rect 10343 24641 10377 24675
rect 10343 24573 10377 24607
rect 10343 24505 10377 24539
rect 10343 24437 10377 24471
rect 10343 24369 10377 24403
rect 10343 24301 10377 24335
rect 10343 24233 10377 24267
rect 10343 24165 10377 24199
rect 10343 24097 10377 24131
rect 10343 24029 10377 24063
rect 10343 23961 10377 23995
rect 10343 23893 10377 23927
rect 10343 23825 10377 23859
rect 23426 23153 23460 23187
rect 23494 23153 23528 23187
rect 23562 23153 23596 23187
rect 23630 23153 23664 23187
rect 23698 23153 23732 23187
rect 23766 23153 23800 23187
rect 34078 23153 34112 23187
rect 34146 23153 34180 23187
rect 34214 23153 34248 23187
rect 34303 23073 34337 23107
rect 34303 23005 34337 23039
rect 34303 22937 34337 22971
rect 34303 22869 34337 22903
rect 34303 22801 34337 22835
rect 34303 22733 34337 22767
rect 34303 22665 34337 22699
rect 34303 22597 34337 22631
rect 34303 22529 34337 22563
rect 34303 22461 34337 22495
rect 34303 22393 34337 22427
rect 34303 22325 34337 22359
rect 34303 22257 34337 22291
rect 34303 22189 34337 22223
rect 34303 22121 34337 22155
rect 34303 22053 34337 22087
rect 34303 21985 34337 22019
rect 34303 21917 34337 21951
rect 34303 21849 34337 21883
rect 34303 21781 34337 21815
rect 34303 21713 34337 21747
rect 34303 21645 34337 21679
rect 34303 21577 34337 21611
rect 34303 21509 34337 21543
rect 34303 21441 34337 21475
rect 34303 21373 34337 21407
rect 34303 21305 34337 21339
rect 34303 21237 34337 21271
rect 34303 21169 34337 21203
rect 34303 21101 34337 21135
rect 34303 21033 34337 21067
rect 34303 20965 34337 20999
rect 34303 20897 34337 20931
rect 34303 20829 34337 20863
rect 34303 20761 34337 20795
rect 34303 20693 34337 20727
rect 34303 20625 34337 20659
rect 34303 20557 34337 20591
rect 34303 20489 34337 20523
rect 34303 20421 34337 20455
rect 34303 20353 34337 20387
rect 34303 20285 34337 20319
rect 34303 20217 34337 20251
rect 34303 20149 34337 20183
rect 34303 20081 34337 20115
rect 34303 20013 34337 20047
rect 34303 19945 34337 19979
rect 34303 19877 34337 19911
rect 34303 19809 34337 19843
rect 34303 19741 34337 19775
rect 34303 19673 34337 19707
rect 34303 19605 34337 19639
rect 34303 19537 34337 19571
rect 34303 19469 34337 19503
rect 34303 19401 34337 19435
rect 34303 19333 34337 19367
rect 34303 19265 34337 19299
rect 34303 19197 34337 19231
rect 34303 19129 34337 19163
rect 34303 19061 34337 19095
rect 34303 18993 34337 19027
rect 34303 18925 34337 18959
rect 34303 18857 34337 18891
rect 34303 18789 34337 18823
rect 34303 18721 34337 18755
rect 34303 18653 34337 18687
rect 34303 18585 34337 18619
rect 34303 18517 34337 18551
rect 34303 18449 34337 18483
rect 34303 18381 34337 18415
rect 34303 18313 34337 18347
rect 34303 18245 34337 18279
rect 34303 18177 34337 18211
rect 34303 18109 34337 18143
rect 34303 18041 34337 18075
rect 34303 17973 34337 18007
rect 34303 17905 34337 17939
rect 34303 17837 34337 17871
rect 34303 17769 34337 17803
rect 34303 17701 34337 17735
rect 34303 17633 34337 17667
rect 34303 17565 34337 17599
rect 34303 17497 34337 17531
rect 34303 17429 34337 17463
rect 34303 17361 34337 17395
rect 34303 17293 34337 17327
rect 34303 17225 34337 17259
rect 34303 17157 34337 17191
rect 34303 17089 34337 17123
rect 34303 17021 34337 17055
rect 34303 16953 34337 16987
rect 34303 16885 34337 16919
rect 34303 16817 34337 16851
rect 34303 16749 34337 16783
rect 34303 16681 34337 16715
rect 34303 16613 34337 16647
rect 23417 16533 23451 16567
rect 23485 16533 23519 16567
rect 23553 16533 23587 16567
rect 23621 16533 23655 16567
rect 23689 16533 23723 16567
rect 23757 16533 23791 16567
rect 23825 16533 23859 16567
rect 23893 16533 23927 16567
rect 23961 16533 23995 16567
rect 24029 16533 24063 16567
rect 24097 16533 24131 16567
rect 24165 16533 24199 16567
rect 24233 16533 24267 16567
rect 24301 16533 24335 16567
rect 24369 16533 24403 16567
rect 24437 16533 24471 16567
rect 24505 16533 24539 16567
rect 24573 16533 24607 16567
rect 24641 16533 24675 16567
rect 24709 16533 24743 16567
rect 24777 16533 24811 16567
rect 24845 16533 24879 16567
rect 24913 16533 24947 16567
rect 24981 16533 25015 16567
rect 25049 16533 25083 16567
rect 25117 16533 25151 16567
rect 25185 16533 25219 16567
rect 25253 16533 25287 16567
rect 25321 16533 25355 16567
rect 25389 16533 25423 16567
rect 25457 16533 25491 16567
rect 25525 16533 25559 16567
rect 25593 16533 25627 16567
rect 25661 16533 25695 16567
rect 25729 16533 25763 16567
rect 25797 16533 25831 16567
rect 25865 16533 25899 16567
rect 25933 16533 25967 16567
rect 26001 16533 26035 16567
rect 26069 16533 26103 16567
rect 26137 16533 26171 16567
rect 26205 16533 26239 16567
rect 26273 16533 26307 16567
rect 26341 16533 26375 16567
rect 26409 16533 26443 16567
rect 26477 16533 26511 16567
rect 26545 16533 26579 16567
rect 26613 16533 26647 16567
rect 26681 16533 26715 16567
rect 26749 16533 26783 16567
rect 26817 16533 26851 16567
rect 26885 16533 26919 16567
rect 26953 16533 26987 16567
rect 27021 16533 27055 16567
rect 27089 16533 27123 16567
rect 27157 16533 27191 16567
rect 27225 16533 27259 16567
rect 27293 16533 27327 16567
rect 27361 16533 27395 16567
rect 27429 16533 27463 16567
rect 27497 16533 27531 16567
rect 27565 16533 27599 16567
rect 27633 16533 27667 16567
rect 27701 16533 27735 16567
rect 27769 16533 27803 16567
rect 27837 16533 27871 16567
rect 27905 16533 27939 16567
rect 27973 16533 28007 16567
rect 28041 16533 28075 16567
rect 28109 16533 28143 16567
rect 28177 16533 28211 16567
rect 28245 16533 28279 16567
rect 28313 16533 28347 16567
rect 28381 16533 28415 16567
rect 28449 16533 28483 16567
rect 28517 16533 28551 16567
rect 28585 16533 28619 16567
rect 28653 16533 28687 16567
rect 28721 16533 28755 16567
rect 28789 16533 28823 16567
rect 28857 16533 28891 16567
rect 28925 16533 28959 16567
rect 28993 16533 29027 16567
rect 29061 16533 29095 16567
rect 29129 16533 29163 16567
rect 29197 16533 29231 16567
rect 29265 16533 29299 16567
rect 29333 16533 29367 16567
rect 29401 16533 29435 16567
rect 29469 16533 29503 16567
rect 29537 16533 29571 16567
rect 29605 16533 29639 16567
rect 29673 16533 29707 16567
rect 29741 16533 29775 16567
rect 29809 16533 29843 16567
rect 29877 16533 29911 16567
rect 29945 16533 29979 16567
rect 30013 16533 30047 16567
rect 30081 16533 30115 16567
rect 30149 16533 30183 16567
rect 30217 16533 30251 16567
rect 30285 16533 30319 16567
rect 30353 16533 30387 16567
rect 30421 16533 30455 16567
rect 30489 16533 30523 16567
rect 30557 16533 30591 16567
rect 30625 16533 30659 16567
rect 30693 16533 30727 16567
rect 30761 16533 30795 16567
rect 30829 16533 30863 16567
rect 30897 16533 30931 16567
rect 30965 16533 30999 16567
rect 31033 16533 31067 16567
rect 31101 16533 31135 16567
rect 31169 16533 31203 16567
rect 31237 16533 31271 16567
rect 31305 16533 31339 16567
rect 31373 16533 31407 16567
rect 31441 16533 31475 16567
rect 31509 16533 31543 16567
rect 31577 16533 31611 16567
rect 31645 16533 31679 16567
rect 31713 16533 31747 16567
rect 31781 16533 31815 16567
rect 31849 16533 31883 16567
rect 31917 16533 31951 16567
rect 31985 16533 32019 16567
rect 32053 16533 32087 16567
rect 32121 16533 32155 16567
rect 32189 16533 32223 16567
rect 32257 16533 32291 16567
rect 32325 16533 32359 16567
rect 32393 16533 32427 16567
rect 32461 16533 32495 16567
rect 32529 16533 32563 16567
rect 32597 16533 32631 16567
rect 32665 16533 32699 16567
rect 32733 16533 32767 16567
rect 32801 16533 32835 16567
rect 32869 16533 32903 16567
rect 32937 16533 32971 16567
rect 33005 16533 33039 16567
rect 33073 16533 33107 16567
rect 33141 16533 33175 16567
rect 33209 16533 33243 16567
rect 33277 16533 33311 16567
rect 33345 16533 33379 16567
rect 33413 16533 33447 16567
rect 33481 16533 33515 16567
rect 33549 16533 33583 16567
rect 33617 16533 33651 16567
rect 33685 16533 33719 16567
rect 33753 16533 33787 16567
rect 33821 16533 33855 16567
rect 33889 16533 33923 16567
rect 33957 16533 33991 16567
rect 34025 16533 34059 16567
rect 34093 16533 34127 16567
rect 34161 16533 34195 16567
rect 34229 16533 34263 16567
rect 5673 13333 5707 13367
rect 5764 13243 5798 13277
rect 5832 13243 5866 13277
rect 5900 13243 5934 13277
rect 5968 13243 6002 13277
rect 6036 13243 6070 13277
rect 6104 13243 6138 13277
rect 6172 13243 6206 13277
rect 6240 13243 6274 13277
rect 6308 13243 6342 13277
rect 6376 13243 6410 13277
rect 6444 13243 6478 13277
rect 6512 13243 6546 13277
rect 6580 13243 6614 13277
rect 6648 13243 6682 13277
rect 6716 13243 6750 13277
rect 6784 13243 6818 13277
rect 6852 13243 6886 13277
rect 6920 13243 6954 13277
rect 6988 13243 7022 13277
rect 7056 13243 7090 13277
rect 7124 13243 7158 13277
rect 7192 13243 7226 13277
rect 7260 13243 7294 13277
rect 7328 13243 7362 13277
rect 7396 13243 7430 13277
rect 7464 13243 7498 13277
rect 7532 13243 7566 13277
rect 7600 13243 7634 13277
rect 7668 13243 7702 13277
rect 7736 13243 7770 13277
rect 7804 13243 7838 13277
rect 7872 13243 7906 13277
rect 7940 13243 7974 13277
rect 8008 13243 8042 13277
rect 8076 13243 8110 13277
rect 8144 13243 8178 13277
rect 8212 13243 8246 13277
rect 8280 13243 8314 13277
rect 8348 13243 8382 13277
rect 8416 13243 8450 13277
rect 8484 13243 8518 13277
rect 8552 13243 8586 13277
rect 8620 13243 8654 13277
rect 8688 13243 8722 13277
rect 8756 13243 8790 13277
rect 8824 13243 8858 13277
rect 8892 13243 8926 13277
rect 8960 13243 8994 13277
rect 9028 13243 9062 13277
rect 9096 13243 9130 13277
rect 9164 13243 9198 13277
rect 9232 13243 9266 13277
rect 9300 13243 9334 13277
rect 9368 13243 9402 13277
rect 9436 13243 9470 13277
rect 9504 13243 9538 13277
rect 9572 13243 9606 13277
rect 9640 13243 9674 13277
rect 9708 13243 9742 13277
rect 9776 13243 9810 13277
rect 9844 13243 9878 13277
rect 9912 13243 9946 13277
rect 9980 13243 10014 13277
rect 10048 13243 10082 13277
rect 10116 13243 10150 13277
rect 10184 13243 10218 13277
rect 10252 13243 10286 13277
<< locali >>
rect 5673 25003 5764 25037
rect 5798 25003 5832 25037
rect 5866 25003 5900 25037
rect 5934 25003 5968 25037
rect 6002 25003 6036 25037
rect 6070 25003 6104 25037
rect 6138 25003 6172 25037
rect 6206 25003 6240 25037
rect 6274 25003 6308 25037
rect 6342 25003 6376 25037
rect 6410 25003 6444 25037
rect 6478 25003 6512 25037
rect 6546 25003 6580 25037
rect 6614 25003 6648 25037
rect 6682 25003 6716 25037
rect 6750 25003 6784 25037
rect 6818 25003 6852 25037
rect 6886 25003 6920 25037
rect 6954 25003 6988 25037
rect 7022 25003 7056 25037
rect 7090 25003 7124 25037
rect 7158 25003 7192 25037
rect 7226 25003 7260 25037
rect 7294 25003 7328 25037
rect 7362 25003 7396 25037
rect 7430 25003 7464 25037
rect 7498 25003 7532 25037
rect 7566 25003 7600 25037
rect 7634 25003 7668 25037
rect 7702 25003 7736 25037
rect 7770 25003 7804 25037
rect 7838 25003 7872 25037
rect 7906 25003 7940 25037
rect 7974 25003 8008 25037
rect 8042 25003 8076 25037
rect 8110 25003 8144 25037
rect 8178 25003 8212 25037
rect 8246 25003 8280 25037
rect 8314 25003 8348 25037
rect 8382 25003 8416 25037
rect 8450 25003 8484 25037
rect 8518 25003 8552 25037
rect 8586 25003 8620 25037
rect 8654 25003 8688 25037
rect 8722 25003 8756 25037
rect 8790 25003 8824 25037
rect 8858 25003 8892 25037
rect 8926 25003 8960 25037
rect 8994 25003 9028 25037
rect 9062 25003 9096 25037
rect 9130 25003 9164 25037
rect 9198 25003 9232 25037
rect 9266 25003 9300 25037
rect 9334 25003 9368 25037
rect 9402 25003 9436 25037
rect 9470 25003 9504 25037
rect 9538 25003 9572 25037
rect 9606 25003 9640 25037
rect 9674 25003 9708 25037
rect 9742 25003 9776 25037
rect 9810 25003 9844 25037
rect 9878 25003 9912 25037
rect 9946 25003 9980 25037
rect 10014 25003 10048 25037
rect 10082 25003 10116 25037
rect 10150 25003 10184 25037
rect 10218 25003 10252 25037
rect 10286 25003 10377 25037
rect 5673 24985 5707 25003
rect 10343 24947 10377 25003
rect 10343 24879 10377 24913
rect 10343 24811 10377 24845
rect 10343 24743 10377 24777
rect 10343 24675 10377 24709
rect 10343 24607 10377 24641
rect 10343 24539 10377 24573
rect 10343 24471 10377 24505
rect 10343 24403 10377 24437
rect 10343 24335 10377 24369
rect 10343 24267 10377 24301
rect 10343 24199 10377 24233
rect 10343 24131 10377 24165
rect 10343 24063 10377 24097
rect 10343 23995 10377 24029
rect 10343 23927 10377 23961
rect 10343 23859 10377 23893
rect 10343 23187 10377 23825
rect 10343 23153 11373 23187
rect 23313 23180 23426 23187
rect 23347 23153 23426 23180
rect 23460 23153 23494 23187
rect 23528 23153 23562 23187
rect 23596 23153 23630 23187
rect 23664 23153 23698 23187
rect 23732 23153 23766 23187
rect 23800 23153 23960 23187
rect 33930 23153 34078 23187
rect 34112 23153 34146 23187
rect 34180 23153 34214 23187
rect 34248 23153 34337 23187
rect 10343 21882 10377 23153
rect 23313 22700 23347 23137
rect 34303 23107 34337 23153
rect 34303 23039 34337 23073
rect 34303 22971 34337 23005
rect 34303 22903 34337 22937
rect 34303 22835 34337 22869
rect 34303 22767 34337 22801
rect 10308 21848 10377 21882
rect 34303 22699 34337 22733
rect 34303 22631 34337 22665
rect 34303 22563 34337 22597
rect 34303 22495 34337 22529
rect 34303 22427 34337 22461
rect 34303 22359 34337 22393
rect 34303 22291 34337 22325
rect 34303 22223 34337 22257
rect 34303 22155 34337 22189
rect 34303 22087 34337 22121
rect 34303 22019 34337 22053
rect 34303 21951 34337 21985
rect 34303 21883 34337 21917
rect 34303 21815 34337 21849
rect 34303 21747 34337 21781
rect 34303 21679 34337 21713
rect 34303 21611 34337 21645
rect 34303 21543 34337 21577
rect 34303 21475 34337 21509
rect 34303 21407 34337 21441
rect 34303 21339 34337 21373
rect 34303 21271 34337 21305
rect 34303 21203 34337 21237
rect 34303 21135 34337 21169
rect 34303 21067 34337 21101
rect 34303 20999 34337 21033
rect 573 20953 658 20987
rect 692 20953 726 20987
rect 760 20953 794 20987
rect 828 20953 862 20987
rect 896 20953 930 20987
rect 964 20953 998 20987
rect 1032 20953 1066 20987
rect 1100 20953 1134 20987
rect 1168 20953 1202 20987
rect 1236 20953 1270 20987
rect 1304 20953 1338 20987
rect 1372 20953 1406 20987
rect 1440 20953 1474 20987
rect 1508 20953 1542 20987
rect 1576 20953 1610 20987
rect 1644 20953 1678 20987
rect 1712 20953 1746 20987
rect 1780 20953 1814 20987
rect 1848 20953 1882 20987
rect 1916 20953 1950 20987
rect 1984 20953 2018 20987
rect 2052 20953 2086 20987
rect 2120 20953 2154 20987
rect 2188 20953 2222 20987
rect 2256 20953 2290 20987
rect 2324 20953 2358 20987
rect 2392 20953 2426 20987
rect 2460 20953 2494 20987
rect 2528 20953 2562 20987
rect 2596 20953 2630 20987
rect 2664 20953 2698 20987
rect 2732 20953 2766 20987
rect 2800 20953 2834 20987
rect 2868 20953 2902 20987
rect 2936 20953 2970 20987
rect 3004 20953 3038 20987
rect 3072 20953 3106 20987
rect 3140 20953 3174 20987
rect 3208 20953 3242 20987
rect 3276 20953 3310 20987
rect 3344 20953 3378 20987
rect 3412 20953 3446 20987
rect 3480 20953 3514 20987
rect 3548 20953 3582 20987
rect 3616 20953 3650 20987
rect 3684 20953 3718 20987
rect 3752 20953 3786 20987
rect 3820 20953 3854 20987
rect 3888 20953 3922 20987
rect 3956 20953 3990 20987
rect 4024 20953 4058 20987
rect 4092 20953 4126 20987
rect 4160 20953 4194 20987
rect 4228 20953 4262 20987
rect 4296 20953 4330 20987
rect 4364 20953 4398 20987
rect 4432 20953 4466 20987
rect 4500 20953 4534 20987
rect 4568 20953 4602 20987
rect 4636 20953 4670 20987
rect 4704 20953 4738 20987
rect 4772 20953 4806 20987
rect 4840 20953 4874 20987
rect 4908 20953 4942 20987
rect 4976 20953 5010 20987
rect 5044 20953 5078 20987
rect 5112 20953 5197 20987
rect 573 20896 607 20953
rect 573 20828 607 20862
rect 573 20760 607 20794
rect 573 20692 607 20726
rect 573 20624 607 20658
rect 573 20556 607 20590
rect 573 20488 607 20522
rect 573 20420 607 20454
rect 573 20352 607 20386
rect 573 20284 607 20318
rect 573 20216 607 20250
rect 573 20148 607 20182
rect 573 20080 607 20114
rect 573 20012 607 20046
rect 573 19944 607 19978
rect 573 19876 607 19910
rect 573 19808 607 19842
rect 573 19740 607 19774
rect 573 19672 607 19706
rect 573 19604 607 19638
rect 573 19536 607 19570
rect 573 19468 607 19502
rect 573 19400 607 19434
rect 573 19332 607 19366
rect 573 19264 607 19298
rect 573 19196 607 19230
rect 573 19128 607 19162
rect 573 19060 607 19094
rect 573 18992 607 19026
rect 573 18924 607 18958
rect 573 18856 607 18890
rect 573 18788 607 18822
rect 573 18720 607 18754
rect 573 18652 607 18686
rect 573 18584 607 18618
rect 573 18516 607 18550
rect 573 18448 607 18482
rect 573 18380 607 18414
rect 573 18312 607 18346
rect 573 18244 607 18278
rect 573 18176 607 18210
rect 573 18108 607 18142
rect 573 18040 607 18074
rect 573 17972 607 18006
rect 573 17904 607 17938
rect 573 17836 607 17870
rect 573 17768 607 17802
rect 573 17700 607 17734
rect 573 17632 607 17666
rect 573 17564 607 17598
rect 573 17496 607 17530
rect 573 17428 607 17462
rect 573 17360 607 17394
rect 573 17292 607 17326
rect 573 17224 607 17258
rect 573 17156 607 17190
rect 573 17088 607 17122
rect 573 17020 607 17054
rect 573 16952 607 16986
rect 573 16884 607 16918
rect 573 16816 607 16850
rect 573 16748 607 16782
rect 573 16680 607 16714
rect 573 16612 607 16646
rect 573 16544 607 16578
rect 573 16476 607 16510
rect 573 16408 607 16442
rect 573 16340 607 16374
rect 573 16272 607 16306
rect 573 16204 607 16238
rect 573 16136 607 16170
rect 573 16068 607 16102
rect 573 16000 607 16034
rect 573 15932 607 15966
rect 573 15864 607 15898
rect 573 15796 607 15830
rect 573 15728 607 15762
rect 573 15660 607 15694
rect 573 15592 607 15626
rect 573 15524 607 15558
rect 573 15456 607 15490
rect 573 15388 607 15422
rect 573 15320 607 15354
rect 573 15252 607 15286
rect 573 15184 607 15218
rect 573 15116 607 15150
rect 573 15048 607 15082
rect 573 14980 607 15014
rect 573 14912 607 14946
rect 573 14844 607 14878
rect 573 14776 607 14810
rect 573 14708 607 14742
rect 573 14640 607 14674
rect 573 14572 607 14606
rect 573 14504 607 14538
rect 573 14436 607 14470
rect 573 14368 607 14402
rect 573 14300 607 14334
rect 573 14232 607 14266
rect 573 14164 607 14198
rect 573 14096 607 14130
rect 573 14028 607 14062
rect 573 13960 607 13994
rect 573 13892 607 13926
rect 573 13824 607 13858
rect 573 13756 607 13790
rect 573 13688 607 13722
rect 573 13620 607 13654
rect 573 13552 607 13586
rect 573 13484 607 13518
rect 573 13416 607 13450
rect 573 13348 607 13382
rect 573 13280 607 13314
rect 573 13212 607 13246
rect 573 13144 607 13178
rect 573 13076 607 13110
rect 573 13008 607 13042
rect 573 12940 607 12974
rect 573 12872 607 12906
rect 573 12804 607 12838
rect 573 12736 607 12770
rect 573 12668 607 12702
rect 573 12600 607 12634
rect 573 12532 607 12566
rect 573 12464 607 12498
rect 573 12396 607 12430
rect 573 12328 607 12362
rect 573 12260 607 12294
rect 573 12192 607 12226
rect 573 12124 607 12158
rect 573 12056 607 12090
rect 573 11988 607 12022
rect 573 11920 607 11954
rect 573 11852 607 11886
rect 573 11784 607 11818
rect 573 11716 607 11750
rect 573 11648 607 11682
rect 573 11557 607 11614
rect 5163 20896 5197 20953
rect 5163 20828 5197 20862
rect 5163 20760 5197 20794
rect 5163 20692 5197 20726
rect 5163 20624 5197 20658
rect 5163 20556 5197 20590
rect 5163 20488 5197 20522
rect 5163 20420 5197 20454
rect 5163 20352 5197 20386
rect 5163 20284 5197 20318
rect 5163 20216 5197 20250
rect 5163 20148 5197 20182
rect 5163 20080 5197 20114
rect 5163 20012 5197 20046
rect 5163 19944 5197 19978
rect 5163 19876 5197 19910
rect 5163 19808 5197 19842
rect 5163 19740 5197 19774
rect 5163 19672 5197 19706
rect 5163 19604 5197 19638
rect 5163 19536 5197 19570
rect 5163 19468 5197 19502
rect 5163 19400 5197 19434
rect 5163 19332 5197 19366
rect 5163 19264 5197 19298
rect 5163 19196 5197 19230
rect 5163 19128 5197 19162
rect 5163 19060 5197 19094
rect 5163 18992 5197 19026
rect 5163 18924 5197 18958
rect 5163 18856 5197 18890
rect 5163 18788 5197 18822
rect 5163 18720 5197 18754
rect 5163 18652 5197 18686
rect 5163 18584 5197 18618
rect 5163 18516 5197 18550
rect 34303 20931 34337 20965
rect 34303 20863 34337 20897
rect 34303 20795 34337 20829
rect 34303 20727 34337 20761
rect 34303 20659 34337 20693
rect 34303 20591 34337 20625
rect 34303 20523 34337 20557
rect 34303 20455 34337 20489
rect 34303 20387 34337 20421
rect 34303 20319 34337 20353
rect 34303 20251 34337 20285
rect 34303 20183 34337 20217
rect 34303 20115 34337 20149
rect 34303 20047 34337 20081
rect 34303 19979 34337 20013
rect 34303 19911 34337 19945
rect 34303 19843 34337 19877
rect 34303 19775 34337 19809
rect 34303 19707 34337 19741
rect 34303 19639 34337 19673
rect 34303 19571 34337 19605
rect 34303 19503 34337 19537
rect 34303 19435 34337 19469
rect 34303 19367 34337 19401
rect 34303 19299 34337 19333
rect 34303 19231 34337 19265
rect 34303 19163 34337 19197
rect 34303 19095 34337 19129
rect 34303 19027 34337 19061
rect 34303 18959 34337 18993
rect 34303 18891 34337 18925
rect 34303 18823 34337 18857
rect 34303 18755 34337 18789
rect 34303 18687 34337 18721
rect 34303 18619 34337 18653
rect 34303 18551 34337 18585
rect 5163 18448 5197 18482
rect 5163 18380 5197 18414
rect 5163 18312 5197 18346
rect 5163 18244 5197 18278
rect 5163 18176 5197 18210
rect 5163 18108 5197 18142
rect 5163 18040 5197 18074
rect 5163 17972 5197 18006
rect 5163 17904 5197 17938
rect 5163 17836 5197 17870
rect 5163 17768 5197 17802
rect 5163 17700 5197 17734
rect 5163 17632 5197 17666
rect 5163 17564 5197 17598
rect 5163 17496 5197 17530
rect 5163 17428 5197 17462
rect 5163 17360 5197 17394
rect 5163 17292 5197 17326
rect 5163 17224 5197 17258
rect 5163 17156 5197 17190
rect 5163 17088 5197 17122
rect 5163 17020 5197 17054
rect 5163 16952 5197 16986
rect 5163 16884 5197 16918
rect 5163 16816 5197 16850
rect 5163 16748 5197 16782
rect 5163 16680 5197 16714
rect 5163 16612 5197 16646
rect 5163 16544 5197 16578
rect 5163 16476 5197 16510
rect 5163 16408 5197 16442
rect 5163 16340 5197 16374
rect 5163 16272 5197 16306
rect 5163 16204 5197 16238
rect 5163 16136 5197 16170
rect 5163 16068 5197 16102
rect 5163 16000 5197 16034
rect 5163 15932 5197 15966
rect 5163 15864 5197 15898
rect 5163 15796 5197 15830
rect 5163 15728 5197 15762
rect 5163 15660 5197 15694
rect 5163 15592 5197 15626
rect 5163 15524 5197 15558
rect 5163 15456 5197 15490
rect 5163 15388 5197 15422
rect 5163 15320 5197 15354
rect 5163 15252 5197 15286
rect 5163 15184 5197 15218
rect 5163 15116 5197 15150
rect 5163 15048 5197 15082
rect 5163 14980 5197 15014
rect 5163 14912 5197 14946
rect 5163 14844 5197 14878
rect 5163 14776 5197 14810
rect 5163 14708 5197 14742
rect 5163 14640 5197 14674
rect 5163 14572 5197 14606
rect 5163 14504 5197 14538
rect 5163 14436 5197 14470
rect 5163 14368 5197 14402
rect 5163 14300 5197 14334
rect 5163 14232 5197 14266
rect 5163 14164 5197 14198
rect 5163 14096 5197 14130
rect 5163 14028 5197 14062
rect 5163 13960 5197 13994
rect 5163 13892 5197 13926
rect 5163 13824 5197 13858
rect 5163 13756 5197 13790
rect 5163 13688 5197 13722
rect 5163 13620 5197 13654
rect 5163 13552 5197 13586
rect 5163 13484 5197 13518
rect 5163 13416 5197 13450
rect 10320 16567 10343 18523
rect 34303 18483 34337 18517
rect 34303 18415 34337 18449
rect 34303 18347 34337 18381
rect 34303 18279 34337 18313
rect 34303 18211 34337 18245
rect 34303 18143 34337 18177
rect 34303 18075 34337 18109
rect 34303 18007 34337 18041
rect 34303 17939 34337 17973
rect 34303 17871 34337 17905
rect 34303 17803 34337 17837
rect 34303 17735 34337 17769
rect 34303 17667 34337 17701
rect 34303 17599 34337 17633
rect 34303 17531 34337 17565
rect 34303 17463 34337 17497
rect 34303 17395 34337 17429
rect 34303 17327 34337 17361
rect 34303 17259 34337 17293
rect 34303 17191 34337 17225
rect 34303 17123 34337 17157
rect 34303 17055 34337 17089
rect 34303 16987 34337 17021
rect 34303 16919 34337 16953
rect 34303 16851 34337 16885
rect 34303 16783 34337 16817
rect 34303 16715 34337 16749
rect 34303 16647 34337 16681
rect 34303 16567 34337 16613
rect 10320 16533 11342 16567
rect 23347 16533 23417 16567
rect 23451 16533 23485 16567
rect 23519 16533 23553 16567
rect 23587 16533 23621 16567
rect 23655 16533 23689 16567
rect 23723 16533 23757 16567
rect 23791 16533 23825 16567
rect 23859 16533 23893 16567
rect 23927 16533 23961 16567
rect 23995 16533 24029 16567
rect 24063 16533 24097 16567
rect 24131 16533 24165 16567
rect 24199 16533 24233 16567
rect 24267 16533 24301 16567
rect 24335 16533 24369 16567
rect 24403 16533 24437 16567
rect 24471 16533 24505 16567
rect 24539 16533 24573 16567
rect 24607 16533 24641 16567
rect 24675 16533 24709 16567
rect 24743 16533 24777 16567
rect 24811 16533 24845 16567
rect 24879 16533 24913 16567
rect 24947 16533 24981 16567
rect 25015 16533 25049 16567
rect 25083 16533 25117 16567
rect 25151 16533 25185 16567
rect 25219 16533 25253 16567
rect 25287 16533 25321 16567
rect 25355 16533 25389 16567
rect 25423 16533 25457 16567
rect 25491 16533 25525 16567
rect 25559 16533 25593 16567
rect 25627 16533 25661 16567
rect 25695 16533 25729 16567
rect 25763 16533 25797 16567
rect 25831 16533 25865 16567
rect 25899 16533 25933 16567
rect 25967 16533 26001 16567
rect 26035 16533 26069 16567
rect 26103 16533 26137 16567
rect 26171 16533 26205 16567
rect 26239 16533 26273 16567
rect 26307 16533 26341 16567
rect 26375 16533 26409 16567
rect 26443 16533 26477 16567
rect 26511 16533 26545 16567
rect 26579 16533 26613 16567
rect 26647 16533 26681 16567
rect 26715 16533 26749 16567
rect 26783 16533 26817 16567
rect 26851 16533 26885 16567
rect 26919 16533 26953 16567
rect 26987 16533 27021 16567
rect 27055 16533 27089 16567
rect 27123 16533 27157 16567
rect 27191 16533 27225 16567
rect 27259 16533 27293 16567
rect 27327 16533 27361 16567
rect 27395 16533 27429 16567
rect 27463 16533 27497 16567
rect 27531 16533 27565 16567
rect 27599 16533 27633 16567
rect 27667 16533 27701 16567
rect 27735 16533 27769 16567
rect 27803 16533 27837 16567
rect 27871 16533 27905 16567
rect 27939 16533 27973 16567
rect 28007 16533 28041 16567
rect 28075 16533 28109 16567
rect 28143 16533 28177 16567
rect 28211 16533 28245 16567
rect 28279 16533 28313 16567
rect 28347 16533 28381 16567
rect 28415 16533 28449 16567
rect 28483 16533 28517 16567
rect 28551 16533 28585 16567
rect 28619 16533 28653 16567
rect 28687 16533 28721 16567
rect 28755 16533 28789 16567
rect 28823 16533 28857 16567
rect 28891 16533 28925 16567
rect 28959 16533 28993 16567
rect 29027 16533 29061 16567
rect 29095 16533 29129 16567
rect 29163 16533 29197 16567
rect 29231 16533 29265 16567
rect 29299 16533 29333 16567
rect 29367 16533 29401 16567
rect 29435 16533 29469 16567
rect 29503 16533 29537 16567
rect 29571 16533 29605 16567
rect 29639 16533 29673 16567
rect 29707 16533 29741 16567
rect 29775 16533 29809 16567
rect 29843 16533 29877 16567
rect 29911 16533 29945 16567
rect 29979 16533 30013 16567
rect 30047 16533 30081 16567
rect 30115 16533 30149 16567
rect 30183 16533 30217 16567
rect 30251 16533 30285 16567
rect 30319 16533 30353 16567
rect 30387 16533 30421 16567
rect 30455 16533 30489 16567
rect 30523 16533 30557 16567
rect 30591 16533 30625 16567
rect 30659 16533 30693 16567
rect 30727 16533 30761 16567
rect 30795 16533 30829 16567
rect 30863 16533 30897 16567
rect 30931 16533 30965 16567
rect 30999 16533 31033 16567
rect 31067 16533 31101 16567
rect 31135 16533 31169 16567
rect 31203 16533 31237 16567
rect 31271 16533 31305 16567
rect 31339 16533 31373 16567
rect 31407 16533 31441 16567
rect 31475 16533 31509 16567
rect 31543 16533 31577 16567
rect 31611 16533 31645 16567
rect 31679 16533 31713 16567
rect 31747 16533 31781 16567
rect 31815 16533 31849 16567
rect 31883 16533 31917 16567
rect 31951 16533 31985 16567
rect 32019 16533 32053 16567
rect 32087 16533 32121 16567
rect 32155 16533 32189 16567
rect 32223 16533 32257 16567
rect 32291 16533 32325 16567
rect 32359 16533 32393 16567
rect 32427 16533 32461 16567
rect 32495 16533 32529 16567
rect 32563 16533 32597 16567
rect 32631 16533 32665 16567
rect 32699 16533 32733 16567
rect 32767 16533 32801 16567
rect 32835 16533 32869 16567
rect 32903 16533 32937 16567
rect 32971 16533 33005 16567
rect 33039 16533 33073 16567
rect 33107 16533 33141 16567
rect 33175 16533 33209 16567
rect 33243 16533 33277 16567
rect 33311 16533 33345 16567
rect 33379 16533 33413 16567
rect 33447 16533 33481 16567
rect 33515 16533 33549 16567
rect 33583 16533 33617 16567
rect 33651 16533 33685 16567
rect 33719 16533 33753 16567
rect 33787 16533 33821 16567
rect 33855 16533 33889 16567
rect 33923 16533 33957 16567
rect 33991 16533 34025 16567
rect 34059 16533 34093 16567
rect 34127 16533 34161 16567
rect 34195 16533 34229 16567
rect 34263 16533 34337 16567
rect 5163 13348 5197 13382
rect 5163 13280 5197 13314
rect 5163 13212 5197 13246
rect 5673 13396 5744 13430
rect 5673 13367 5707 13396
rect 5673 13277 5707 13333
rect 10320 13330 10343 16533
rect 34580 16447 34710 16530
rect 34580 16413 34623 16447
rect 34657 16413 34710 16447
rect 34580 16400 34710 16413
rect 10310 13277 10343 13330
rect 5673 13243 5764 13277
rect 5798 13243 5832 13277
rect 5866 13243 5900 13277
rect 5934 13243 5968 13277
rect 6002 13243 6036 13277
rect 6070 13243 6104 13277
rect 6138 13243 6172 13277
rect 6206 13243 6240 13277
rect 6274 13243 6308 13277
rect 6342 13243 6376 13277
rect 6410 13243 6444 13277
rect 6478 13243 6512 13277
rect 6546 13243 6580 13277
rect 6614 13243 6648 13277
rect 6682 13243 6716 13277
rect 6750 13243 6784 13277
rect 6818 13243 6852 13277
rect 6886 13243 6920 13277
rect 6954 13243 6988 13277
rect 7022 13243 7056 13277
rect 7090 13243 7124 13277
rect 7158 13243 7192 13277
rect 7226 13243 7260 13277
rect 7294 13243 7328 13277
rect 7362 13243 7396 13277
rect 7430 13243 7464 13277
rect 7498 13243 7532 13277
rect 7566 13243 7600 13277
rect 7634 13243 7668 13277
rect 7702 13243 7736 13277
rect 7770 13243 7804 13277
rect 7838 13243 7872 13277
rect 7906 13243 7940 13277
rect 7974 13243 8008 13277
rect 8042 13243 8076 13277
rect 8110 13243 8144 13277
rect 8178 13243 8212 13277
rect 8246 13243 8280 13277
rect 8314 13243 8348 13277
rect 8382 13243 8416 13277
rect 8450 13243 8484 13277
rect 8518 13243 8552 13277
rect 8586 13243 8620 13277
rect 8654 13243 8688 13277
rect 8722 13243 8756 13277
rect 8790 13243 8824 13277
rect 8858 13243 8892 13277
rect 8926 13243 8960 13277
rect 8994 13243 9028 13277
rect 9062 13243 9096 13277
rect 9130 13243 9164 13277
rect 9198 13243 9232 13277
rect 9266 13243 9300 13277
rect 9334 13243 9368 13277
rect 9402 13243 9436 13277
rect 9470 13243 9504 13277
rect 9538 13243 9572 13277
rect 9606 13243 9640 13277
rect 9674 13243 9708 13277
rect 9742 13243 9776 13277
rect 9810 13243 9844 13277
rect 9878 13243 9912 13277
rect 9946 13243 9980 13277
rect 10014 13243 10048 13277
rect 10082 13243 10116 13277
rect 10150 13243 10184 13277
rect 10218 13243 10252 13277
rect 10286 13243 10343 13277
rect 5163 13144 5197 13178
rect 5163 13076 5197 13110
rect 5163 13008 5197 13042
rect 5163 12940 5197 12974
rect 5163 12872 5197 12906
rect 5163 12804 5197 12838
rect 5163 12736 5197 12770
rect 5163 12668 5197 12702
rect 5163 12600 5197 12634
rect 5163 12532 5197 12566
rect 5163 12464 5197 12498
rect 5163 12396 5197 12430
rect 5163 12328 5197 12362
rect 5163 12260 5197 12294
rect 5163 12192 5197 12226
rect 5163 12124 5197 12158
rect 5163 12056 5197 12090
rect 5163 11988 5197 12022
rect 5163 11920 5197 11954
rect 5163 11852 5197 11886
rect 5163 11784 5197 11818
rect 5163 11716 5197 11750
rect 5163 11648 5197 11682
rect 5163 11557 5197 11614
rect 573 11523 658 11557
rect 692 11523 726 11557
rect 760 11523 794 11557
rect 828 11523 862 11557
rect 896 11523 930 11557
rect 964 11523 998 11557
rect 1032 11523 1066 11557
rect 1100 11523 1134 11557
rect 1168 11523 1202 11557
rect 1236 11523 1270 11557
rect 1304 11523 1338 11557
rect 1372 11523 1406 11557
rect 1440 11523 1474 11557
rect 1508 11523 1542 11557
rect 1576 11523 1610 11557
rect 1644 11523 1678 11557
rect 1712 11523 1746 11557
rect 1780 11523 1814 11557
rect 1848 11523 1882 11557
rect 1916 11523 1950 11557
rect 1984 11523 2018 11557
rect 2052 11523 2086 11557
rect 2120 11523 2154 11557
rect 2188 11523 2222 11557
rect 2256 11523 2290 11557
rect 2324 11523 2358 11557
rect 2392 11523 2426 11557
rect 2460 11523 2494 11557
rect 2528 11523 2562 11557
rect 2596 11523 2630 11557
rect 2664 11523 2698 11557
rect 2732 11523 2766 11557
rect 2800 11523 2834 11557
rect 2868 11523 2902 11557
rect 2936 11523 2970 11557
rect 3004 11523 3038 11557
rect 3072 11523 3106 11557
rect 3140 11523 3174 11557
rect 3208 11523 3242 11557
rect 3276 11523 3310 11557
rect 3344 11523 3378 11557
rect 3412 11523 3446 11557
rect 3480 11523 3514 11557
rect 3548 11523 3582 11557
rect 3616 11523 3650 11557
rect 3684 11523 3718 11557
rect 3752 11523 3786 11557
rect 3820 11523 3854 11557
rect 3888 11523 3922 11557
rect 3956 11523 3990 11557
rect 4024 11523 4058 11557
rect 4092 11523 4126 11557
rect 4160 11523 4194 11557
rect 4228 11523 4262 11557
rect 4296 11523 4330 11557
rect 4364 11523 4398 11557
rect 4432 11523 4466 11557
rect 4500 11523 4534 11557
rect 4568 11523 4602 11557
rect 4636 11523 4670 11557
rect 4704 11523 4738 11557
rect 4772 11523 4806 11557
rect 4840 11523 4874 11557
rect 4908 11523 4942 11557
rect 4976 11523 5010 11557
rect 5044 11523 5078 11557
rect 5112 11523 5197 11557
<< viali >>
rect 34623 16413 34657 16447
<< metal1 >>
rect 10340 17650 10343 17720
rect 34580 16447 34710 16480
rect 34580 16413 34623 16447
rect 34657 16413 34710 16447
rect 34580 16400 34710 16413
rect 34580 15220 34640 16400
rect 34580 15156 34680 15220
rect 34580 15104 34604 15156
rect 34656 15104 34680 15156
rect 34580 15011 34680 15104
rect 34580 14959 34604 15011
rect 34656 14959 34680 15011
rect 34580 14920 34680 14959
rect 17100 7740 17110 7770
rect 14780 6656 15078 7438
rect 15940 6660 16240 7440
rect 17100 6660 17400 7740
<< via1 >>
rect 34604 15104 34656 15156
rect 34604 14959 34656 15011
<< metal2 >>
rect 34580 15158 34680 15220
rect 34580 15102 34602 15158
rect 34658 15102 34680 15158
rect 34580 15013 34680 15102
rect 34580 14957 34602 15013
rect 34658 14957 34680 15013
rect 34580 14920 34680 14957
rect 5673 13396 5744 13430
rect 4080 12200 4384 12260
rect 4090 12080 4394 12140
<< via2 >>
rect 34602 15156 34658 15158
rect 34602 15104 34604 15156
rect 34604 15104 34656 15156
rect 34656 15104 34658 15156
rect 34602 15102 34658 15104
rect 34602 15011 34658 15013
rect 34602 14959 34604 15011
rect 34604 14959 34656 15011
rect 34656 14959 34658 15011
rect 34602 14957 34658 14959
<< metal3 >>
rect 34580 15162 34680 15220
rect 34580 15098 34598 15162
rect 34662 15098 34680 15162
rect 34580 15017 34680 15098
rect 34580 14953 34598 15017
rect 34662 14953 34680 15017
rect 34580 14920 34680 14953
<< via3 >>
rect 34598 15158 34662 15162
rect 34598 15102 34602 15158
rect 34602 15102 34658 15158
rect 34658 15102 34662 15158
rect 34598 15098 34662 15102
rect 34598 15013 34662 15017
rect 34598 14957 34602 15013
rect 34602 14957 34658 15013
rect 34658 14957 34662 15013
rect 34598 14953 34662 14957
<< metal4 >>
rect 0 25220 300 25520
rect 40880 16150 41180 16450
rect 40890 15890 41560 16070
rect 41260 15770 41560 15890
rect 34590 15162 34670 15180
rect 34590 15098 34598 15162
rect 34662 15098 34670 15162
rect 34590 15080 34670 15098
rect 34590 15017 34670 15030
rect 34590 14953 34598 15017
rect 34662 14953 34670 15017
rect 34590 14940 34670 14953
rect 33640 13910 33680 14010
rect 120 11180 420 11480
rect 10010 10840 10310 11140
rect 10010 10350 10310 10650
rect 4320 880 4620 1180
rect 4820 880 5120 1180
rect 10120 330 10420 630
rect 33140 -30 33440 270
use 2stage_op_amp  2stage_op_amp_1
timestamp 1757161594
transform 1 0 10950 0 1 140
box -11080 -340 30862 25583
<< labels >>
flabel metal4 s 120 11180 420 11480 0 FreeSans 1562 0 0 0 Rgm
port 1 nsew
flabel metal4 s 40880 16150 41180 16450 0 FreeSans 1562 0 0 0 Vop
port 2 nsew
flabel metal4 s 10010 10840 10310 11140 0 FreeSans 1562 0 0 0 Vm
port 3 nsew
flabel metal4 s 4320 880 4620 1180 0 FreeSans 1562 0 0 0 en_1
port 4 nsew
flabel metal4 s 0 25220 300 25520 0 FreeSans 1562 0 0 0 Vdd
port 5 nsew
flabel metal4 s 10120 330 10420 630 0 FreeSans 1562 0 0 0 Vss
port 6 nsew
flabel metal4 s 33140 -30 33440 270 0 FreeSans 1562 0 0 0 Vref
port 7 nsew
flabel metal4 s 4820 880 5120 1180 0 FreeSans 1562 0 0 0 en_2
port 8 nsew
flabel metal4 s 41260 15770 41560 16070 0 FreeSans 1562 0 0 0 Vom
port 9 nsew
flabel metal4 s 10010 10350 10310 10650 0 FreeSans 1562 0 0 0 Vp
port 10 nsew
<< end >>
