magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -184 -257 184 195
<< nmoslvt >>
rect -100 -231 100 169
<< ndiff >>
rect -158 88 -100 169
rect -158 54 -146 88
rect -112 54 -100 88
rect -158 20 -100 54
rect -158 -14 -146 20
rect -112 -14 -100 20
rect -158 -48 -100 -14
rect -158 -82 -146 -48
rect -112 -82 -100 -48
rect -158 -116 -100 -82
rect -158 -150 -146 -116
rect -112 -150 -100 -116
rect -158 -231 -100 -150
rect 100 88 158 169
rect 100 54 112 88
rect 146 54 158 88
rect 100 20 158 54
rect 100 -14 112 20
rect 146 -14 158 20
rect 100 -48 158 -14
rect 100 -82 112 -48
rect 146 -82 158 -48
rect 100 -116 158 -82
rect 100 -150 112 -116
rect 146 -150 158 -116
rect 100 -231 158 -150
<< ndiffc >>
rect -146 54 -112 88
rect -146 -14 -112 20
rect -146 -82 -112 -48
rect -146 -150 -112 -116
rect 112 54 146 88
rect 112 -14 146 20
rect 112 -82 146 -48
rect 112 -150 146 -116
<< poly >>
rect -75 241 75 257
rect -75 224 -51 241
rect -100 207 -51 224
rect -17 207 17 241
rect 51 224 75 241
rect 51 207 100 224
rect -100 169 100 207
rect -100 -257 100 -231
<< polycont >>
rect -51 207 -17 241
rect 17 207 51 241
<< locali >>
rect -75 207 -53 241
rect -17 207 17 241
rect 53 207 75 241
rect -146 94 -112 117
rect -146 22 -112 54
rect -146 -48 -112 -14
rect -146 -116 -112 -84
rect -146 -179 -112 -156
rect 112 94 146 117
rect 112 22 146 54
rect 112 -48 146 -14
rect 112 -116 146 -84
rect 112 -179 146 -156
<< viali >>
rect -53 207 -51 241
rect -51 207 -19 241
rect 19 207 51 241
rect 51 207 53 241
rect -146 88 -112 94
rect -146 60 -112 88
rect -146 20 -112 22
rect -146 -12 -112 20
rect -146 -82 -112 -50
rect -146 -84 -112 -82
rect -146 -150 -112 -122
rect -146 -156 -112 -150
rect 112 88 146 94
rect 112 60 146 88
rect 112 20 146 22
rect 112 -12 146 20
rect 112 -82 146 -50
rect 112 -84 146 -82
rect 112 -150 146 -122
rect 112 -156 146 -150
<< metal1 >>
rect -71 241 71 247
rect -71 207 -53 241
rect -19 207 19 241
rect 53 207 71 241
rect -71 201 71 207
rect -152 94 -106 113
rect -152 60 -146 94
rect -112 60 -106 94
rect -152 22 -106 60
rect -152 -12 -146 22
rect -112 -12 -106 22
rect -152 -50 -106 -12
rect -152 -84 -146 -50
rect -112 -84 -106 -50
rect -152 -122 -106 -84
rect -152 -156 -146 -122
rect -112 -156 -106 -122
rect -152 -175 -106 -156
rect 106 94 152 113
rect 106 60 112 94
rect 146 60 152 94
rect 106 22 152 60
rect 106 -12 112 22
rect 146 -12 152 22
rect 106 -50 152 -12
rect 106 -84 112 -50
rect 146 -84 152 -50
rect 106 -122 152 -84
rect 106 -156 112 -122
rect 146 -156 152 -122
rect 106 -175 152 -156
<< end >>
