magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -726 4504 1246 4596
rect -726 -304 -634 4504
rect 1154 -304 1246 4504
rect -726 -436 1246 -304
<< psubdiff >>
rect -700 4530 1220 4570
rect -700 -330 -660 4530
rect 1180 -330 1220 4530
rect -700 -353 1220 -330
rect -700 -387 -641 -353
rect -607 -387 -573 -353
rect -539 -387 -505 -353
rect -471 -387 -437 -353
rect -403 -387 -369 -353
rect -335 -387 -301 -353
rect -267 -387 -233 -353
rect -199 -387 -165 -353
rect -131 -387 -97 -353
rect -63 -387 -29 -353
rect 5 -387 39 -353
rect 73 -387 107 -353
rect 141 -387 175 -353
rect 209 -387 243 -353
rect 277 -387 311 -353
rect 345 -387 379 -353
rect 413 -387 447 -353
rect 481 -387 515 -353
rect 549 -387 583 -353
rect 617 -387 651 -353
rect 685 -387 719 -353
rect 753 -387 787 -353
rect 821 -387 855 -353
rect 889 -387 923 -353
rect 957 -387 991 -353
rect 1025 -387 1059 -353
rect 1093 -387 1127 -353
rect 1161 -387 1220 -353
rect -700 -410 1220 -387
<< psubdiffcont >>
rect -641 -387 -607 -353
rect -573 -387 -539 -353
rect -505 -387 -471 -353
rect -437 -387 -403 -353
rect -369 -387 -335 -353
rect -301 -387 -267 -353
rect -233 -387 -199 -353
rect -165 -387 -131 -353
rect -97 -387 -63 -353
rect -29 -387 5 -353
rect 39 -387 73 -353
rect 107 -387 141 -353
rect 175 -387 209 -353
rect 243 -387 277 -353
rect 311 -387 345 -353
rect 379 -387 413 -353
rect 447 -387 481 -353
rect 515 -387 549 -353
rect 583 -387 617 -353
rect 651 -387 685 -353
rect 719 -387 753 -353
rect 787 -387 821 -353
rect 855 -387 889 -353
rect 923 -387 957 -353
rect 991 -387 1025 -353
rect 1059 -387 1093 -353
rect 1127 -387 1161 -353
<< locali >>
rect -700 4530 1220 4570
rect -700 -330 -660 4530
rect 1180 -330 1220 4530
rect -700 -353 1220 -330
rect -700 -387 -657 -353
rect -607 -387 -585 -353
rect -539 -387 -513 -353
rect -471 -387 -441 -353
rect -403 -387 -369 -353
rect -335 -387 -301 -353
rect -263 -387 -233 -353
rect -191 -387 -165 -353
rect -119 -387 -97 -353
rect -47 -387 -29 -353
rect 25 -387 39 -353
rect 97 -387 107 -353
rect 169 -387 175 -353
rect 241 -387 243 -353
rect 277 -387 279 -353
rect 345 -387 351 -353
rect 413 -387 423 -353
rect 481 -387 495 -353
rect 549 -387 567 -353
rect 617 -387 639 -353
rect 685 -387 711 -353
rect 753 -387 783 -353
rect 821 -387 855 -353
rect 889 -387 923 -353
rect 961 -387 991 -353
rect 1033 -387 1059 -353
rect 1105 -387 1127 -353
rect 1177 -387 1220 -353
rect -700 -410 1220 -387
<< viali >>
rect -657 -387 -641 -353
rect -641 -387 -623 -353
rect -585 -387 -573 -353
rect -573 -387 -551 -353
rect -513 -387 -505 -353
rect -505 -387 -479 -353
rect -441 -387 -437 -353
rect -437 -387 -407 -353
rect -369 -387 -335 -353
rect -297 -387 -267 -353
rect -267 -387 -263 -353
rect -225 -387 -199 -353
rect -199 -387 -191 -353
rect -153 -387 -131 -353
rect -131 -387 -119 -353
rect -81 -387 -63 -353
rect -63 -387 -47 -353
rect -9 -387 5 -353
rect 5 -387 25 -353
rect 63 -387 73 -353
rect 73 -387 97 -353
rect 135 -387 141 -353
rect 141 -387 169 -353
rect 207 -387 209 -353
rect 209 -387 241 -353
rect 279 -387 311 -353
rect 311 -387 313 -353
rect 351 -387 379 -353
rect 379 -387 385 -353
rect 423 -387 447 -353
rect 447 -387 457 -353
rect 495 -387 515 -353
rect 515 -387 529 -353
rect 567 -387 583 -353
rect 583 -387 601 -353
rect 639 -387 651 -353
rect 651 -387 673 -353
rect 711 -387 719 -353
rect 719 -387 745 -353
rect 783 -387 787 -353
rect 787 -387 817 -353
rect 855 -387 889 -353
rect 927 -387 957 -353
rect 957 -387 961 -353
rect 999 -387 1025 -353
rect 1025 -387 1033 -353
rect 1071 -387 1093 -353
rect 1093 -387 1105 -353
rect 1143 -387 1161 -353
rect 1161 -387 1177 -353
<< metal1 >>
rect -580 4420 1120 4480
rect -460 4320 -380 4420
rect -160 4320 -80 4420
rect 140 4320 220 4420
rect 440 4320 520 4420
rect 740 4320 820 4420
rect 1040 4320 1120 4420
rect -580 4260 -380 4320
rect -260 4260 -80 4320
rect 20 4260 220 4320
rect 320 4260 520 4320
rect 620 4260 820 4320
rect 920 4260 1120 4320
rect -140 4224 -60 4229
rect -144 4220 -59 4224
rect -144 4168 -128 4220
rect -76 4168 -59 4220
rect -144 4165 -59 4168
rect 157 4220 242 4224
rect 157 4168 173 4220
rect 225 4168 242 4220
rect 157 4165 242 4168
rect 456 4218 541 4222
rect 456 4166 472 4218
rect 524 4166 541 4218
rect 756 4221 841 4225
rect 756 4169 772 4221
rect 824 4169 841 4221
rect 756 4166 841 4169
rect -560 4060 -380 4120
rect -288 4119 -175 4121
rect -288 4067 -258 4119
rect -206 4067 -175 4119
rect -288 4065 -175 4067
rect -460 4040 -380 4060
rect -440 80 -380 4040
rect -140 100 -60 4165
rect 160 4120 240 4165
rect 456 4163 541 4166
rect 460 4120 540 4163
rect 20 4060 240 4120
rect 320 4060 540 4120
rect 613 4118 726 4120
rect 613 4066 643 4118
rect 695 4066 726 4118
rect 613 4064 726 4066
rect 140 4020 240 4060
rect 440 4040 540 4060
rect 160 100 240 4020
rect 460 100 540 4040
rect 760 100 840 4166
rect 1040 4120 1120 4260
rect 920 4060 1120 4120
rect 1040 4040 1120 4060
rect 1060 80 1120 4040
rect -460 60 -380 80
rect 1040 60 1120 80
rect -560 48 -380 60
rect -565 44 -380 48
rect -565 -8 -549 44
rect -497 0 -380 44
rect -263 40 -178 42
rect -280 38 -178 40
rect 40 38 120 40
rect -497 -8 -480 0
rect -565 -11 -480 -8
rect -560 -50 -480 -11
rect -280 -14 -247 38
rect -195 -14 -178 38
rect -280 -17 -178 -14
rect 32 34 120 38
rect 340 36 420 40
rect 640 39 720 40
rect -280 -50 -180 -17
rect 32 -18 48 34
rect 100 -18 120 34
rect 32 -21 120 -18
rect 40 -50 120 -21
rect 335 32 420 36
rect 335 -20 351 32
rect 403 -20 420 32
rect 634 35 720 39
rect 940 37 1120 60
rect 634 -17 650 35
rect 702 -17 720 35
rect 634 -20 720 -17
rect 335 -23 420 -20
rect 340 -50 420 -23
rect 640 -50 720 -20
rect 932 33 1120 37
rect 932 -19 948 33
rect 1000 0 1120 33
rect 1000 -19 1020 0
rect 932 -22 1020 -19
rect 940 -50 1020 -22
rect -560 -110 -380 -50
rect -280 -110 -80 -50
rect 20 -110 220 -50
rect 340 -110 520 -50
rect 640 -110 820 -50
rect 920 -110 1120 -50
rect -460 -210 -380 -110
rect -160 -210 -80 -110
rect 140 -210 220 -110
rect 440 -210 520 -110
rect 740 -210 820 -110
rect 1040 -210 1120 -110
rect -580 -270 -380 -210
rect -280 -270 -80 -210
rect 20 -270 220 -210
rect 340 -270 520 -210
rect 640 -270 820 -210
rect 920 -270 1120 -210
rect -700 -353 1220 -330
rect -700 -387 -657 -353
rect -623 -387 -585 -353
rect -551 -387 -513 -353
rect -479 -387 -441 -353
rect -407 -387 -369 -353
rect -335 -387 -297 -353
rect -263 -387 -225 -353
rect -191 -387 -153 -353
rect -119 -387 -81 -353
rect -47 -387 -9 -353
rect 25 -387 63 -353
rect 97 -387 135 -353
rect 169 -387 207 -353
rect 241 -387 279 -353
rect 313 -387 351 -353
rect 385 -387 423 -353
rect 457 -387 495 -353
rect 529 -387 567 -353
rect 601 -387 639 -353
rect 673 -387 711 -353
rect 745 -387 783 -353
rect 817 -387 855 -353
rect 889 -387 927 -353
rect 961 -387 999 -353
rect 1033 -387 1071 -353
rect 1105 -387 1143 -353
rect 1177 -387 1220 -353
rect -700 -410 1220 -387
<< via1 >>
rect -128 4168 -76 4220
rect 173 4168 225 4220
rect 472 4166 524 4218
rect 772 4169 824 4221
rect -258 4067 -206 4119
rect 643 4066 695 4118
rect -549 -8 -497 44
rect -247 -14 -195 38
rect 48 -18 100 34
rect 351 -20 403 32
rect 650 -17 702 35
rect 948 -19 1000 33
<< metal2 >>
rect -790 4230 -700 4240
rect -134 4230 -69 4234
rect 167 4230 232 4234
rect 466 4230 531 4232
rect 766 4230 831 4235
rect -790 4221 840 4230
rect -790 4220 772 4221
rect -790 4168 -128 4220
rect -76 4168 173 4220
rect 225 4218 772 4220
rect 225 4168 472 4218
rect -790 4166 472 4168
rect 524 4169 772 4218
rect 824 4169 840 4221
rect 524 4166 840 4169
rect -790 4160 840 4166
rect -278 4130 -185 4131
rect -700 4119 720 4130
rect -700 4067 -258 4119
rect -206 4118 720 4119
rect -206 4067 643 4118
rect -700 4066 643 4067
rect 695 4066 720 4118
rect -700 4060 720 4066
rect -278 4055 -185 4060
rect 623 4054 716 4060
rect -555 44 -490 58
rect -555 40 -549 44
rect -580 -8 -549 40
rect -497 40 -490 44
rect -253 40 -188 52
rect 42 40 107 48
rect 345 40 410 46
rect 644 40 709 49
rect 942 40 1007 47
rect -497 38 1020 40
rect -497 -8 -247 38
rect -580 -14 -247 -8
rect -195 35 1020 38
rect -195 34 650 35
rect -195 -14 48 34
rect -580 -18 48 -14
rect 100 32 650 34
rect 100 -18 351 32
rect -580 -20 351 -18
rect 403 -17 650 32
rect 702 33 1020 35
rect 702 -17 948 33
rect 403 -19 948 -17
rect 1000 -19 1020 33
rect 403 -20 1020 -19
rect -580 -40 1020 -20
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_0
timestamp 1757161594
transform 0 1 107 -1 0 4368
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_1
timestamp 1757161594
transform 0 1 -193 -1 0 -162
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_2
timestamp 1757161594
transform 0 1 107 -1 0 -162
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_3
timestamp 1757161594
transform 0 1 407 -1 0 -162
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_4
timestamp 1757161594
transform 0 1 707 -1 0 -162
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_5
timestamp 1757161594
transform 0 1 -193 -1 0 4368
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_6
timestamp 1757161594
transform 0 1 407 -1 0 4368
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_7
timestamp 1757161594
transform 0 1 707 -1 0 4368
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_8
timestamp 1757161594
transform 0 1 1007 -1 0 -162
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_9
timestamp 1757161594
transform 0 1 1007 -1 0 4368
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_10
timestamp 1757161594
transform 0 1 -493 -1 0 -162
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_BX6RT7  sky130_fd_pr__nfet_01v8_lvt_BX6RT7_11
timestamp 1757161594
transform 0 1 -493 -1 0 4368
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_N42WW9  sky130_fd_pr__nfet_01v8_lvt_N42WW9_0
timestamp 1757161594
transform 0 1 -193 -1 0 2058
box -2084 -107 2084 107
use sky130_fd_pr__nfet_01v8_lvt_N42WW9  sky130_fd_pr__nfet_01v8_lvt_N42WW9_1
timestamp 1757161594
transform 0 1 107 -1 0 2058
box -2084 -107 2084 107
use sky130_fd_pr__nfet_01v8_lvt_N42WW9  sky130_fd_pr__nfet_01v8_lvt_N42WW9_2
timestamp 1757161594
transform 0 1 407 -1 0 2058
box -2084 -107 2084 107
use sky130_fd_pr__nfet_01v8_lvt_N42WW9  sky130_fd_pr__nfet_01v8_lvt_N42WW9_3
timestamp 1757161594
transform 0 1 707 -1 0 2058
box -2084 -107 2084 107
use sky130_fd_pr__nfet_01v8_lvt_N42WW9  sky130_fd_pr__nfet_01v8_lvt_N42WW9_4
timestamp 1757161594
transform 0 1 1007 -1 0 2058
box -2084 -107 2084 107
use sky130_fd_pr__nfet_01v8_lvt_N42WW9  sky130_fd_pr__nfet_01v8_lvt_N42WW9_5
timestamp 1757161594
transform 0 1 -493 -1 0 2058
box -2084 -107 2084 107
<< end >>
