magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< error_p >>
rect -36 145 36 151
rect -36 111 -17 145
rect -36 105 36 111
<< nwell >>
rect -144 -198 144 164
<< pmoslvt >>
rect -50 -136 50 64
<< pdiff >>
rect -108 15 -50 64
rect -108 -19 -96 15
rect -62 -19 -50 15
rect -108 -53 -50 -19
rect -108 -87 -96 -53
rect -62 -87 -50 -53
rect -108 -136 -50 -87
rect 50 15 108 64
rect 50 -19 62 15
rect 96 -19 108 15
rect 50 -53 108 -19
rect 50 -87 62 -53
rect 96 -87 108 -53
rect 50 -136 108 -87
<< pdiffc >>
rect -96 -19 -62 15
rect -96 -87 -62 -53
rect 62 -19 96 15
rect 62 -87 96 -53
<< poly >>
rect -40 145 40 161
rect -40 128 -17 145
rect -50 111 -17 128
rect 17 128 40 145
rect 17 111 50 128
rect -50 64 50 111
rect -50 -162 50 -136
<< polycont >>
rect -17 111 17 145
<< locali >>
rect -40 111 -17 145
rect 17 111 40 145
rect -96 17 -62 42
rect -96 -53 -62 -19
rect -96 -114 -62 -89
rect 62 17 96 42
rect 62 -53 96 -19
rect 62 -114 96 -89
<< viali >>
rect -17 111 17 145
rect -96 15 -62 17
rect -96 -17 -62 15
rect -96 -87 -62 -55
rect -96 -89 -62 -87
rect 62 15 96 17
rect 62 -17 96 15
rect 62 -87 96 -55
rect 62 -89 96 -87
<< metal1 >>
rect -36 145 36 151
rect -36 111 -17 145
rect 17 111 36 145
rect -36 105 36 111
rect -102 17 -56 38
rect -102 -17 -96 17
rect -62 -17 -56 17
rect -102 -55 -56 -17
rect -102 -89 -96 -55
rect -62 -89 -56 -55
rect -102 -110 -56 -89
rect 56 17 102 38
rect 56 -17 62 17
rect 96 -17 102 17
rect 56 -55 102 -17
rect 56 -89 62 -55
rect 96 -89 102 -55
rect 56 -110 102 -89
<< end >>
