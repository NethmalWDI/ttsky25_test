magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -1084 -107 1084 45
<< nmoslvt >>
rect -1000 -81 1000 19
<< ndiff >>
rect -1058 -14 -1000 19
rect -1058 -48 -1046 -14
rect -1012 -48 -1000 -14
rect -1058 -81 -1000 -48
rect 1000 -14 1058 19
rect 1000 -48 1012 -14
rect 1046 -48 1058 -14
rect 1000 -81 1058 -48
<< ndiffc >>
rect -1046 -48 -1012 -14
rect 1012 -48 1046 -14
<< poly >>
rect -705 91 705 107
rect -705 74 -663 91
rect -1000 57 -663 74
rect -629 57 -595 91
rect -561 57 -527 91
rect -493 57 -459 91
rect -425 57 -391 91
rect -357 57 -323 91
rect -289 57 -255 91
rect -221 57 -187 91
rect -153 57 -119 91
rect -85 57 -51 91
rect -17 57 17 91
rect 51 57 85 91
rect 119 57 153 91
rect 187 57 221 91
rect 255 57 289 91
rect 323 57 357 91
rect 391 57 425 91
rect 459 57 493 91
rect 527 57 561 91
rect 595 57 629 91
rect 663 74 705 91
rect 663 57 1000 74
rect -1000 19 1000 57
rect -1000 -107 1000 -81
<< polycont >>
rect -663 57 -629 91
rect -595 57 -561 91
rect -527 57 -493 91
rect -459 57 -425 91
rect -391 57 -357 91
rect -323 57 -289 91
rect -255 57 -221 91
rect -187 57 -153 91
rect -119 57 -85 91
rect -51 57 -17 91
rect 17 57 51 91
rect 85 57 119 91
rect 153 57 187 91
rect 221 57 255 91
rect 289 57 323 91
rect 357 57 391 91
rect 425 57 459 91
rect 493 57 527 91
rect 561 57 595 91
rect 629 57 663 91
<< locali >>
rect -705 57 -665 91
rect -629 57 -595 91
rect -559 57 -527 91
rect -487 57 -459 91
rect -415 57 -391 91
rect -343 57 -323 91
rect -271 57 -255 91
rect -199 57 -187 91
rect -127 57 -119 91
rect -55 57 -51 91
rect 51 57 55 91
rect 119 57 127 91
rect 187 57 199 91
rect 255 57 271 91
rect 323 57 343 91
rect 391 57 415 91
rect 459 57 487 91
rect 527 57 559 91
rect 595 57 629 91
rect 665 57 705 91
rect -1046 -14 -1012 12
rect -1046 -74 -1012 -48
rect 1012 -14 1046 12
rect 1012 -74 1046 -48
<< viali >>
rect -665 57 -663 91
rect -663 57 -631 91
rect -593 57 -561 91
rect -561 57 -559 91
rect -521 57 -493 91
rect -493 57 -487 91
rect -449 57 -425 91
rect -425 57 -415 91
rect -377 57 -357 91
rect -357 57 -343 91
rect -305 57 -289 91
rect -289 57 -271 91
rect -233 57 -221 91
rect -221 57 -199 91
rect -161 57 -153 91
rect -153 57 -127 91
rect -89 57 -85 91
rect -85 57 -55 91
rect -17 57 17 91
rect 55 57 85 91
rect 85 57 89 91
rect 127 57 153 91
rect 153 57 161 91
rect 199 57 221 91
rect 221 57 233 91
rect 271 57 289 91
rect 289 57 305 91
rect 343 57 357 91
rect 357 57 377 91
rect 415 57 425 91
rect 425 57 449 91
rect 487 57 493 91
rect 493 57 521 91
rect 559 57 561 91
rect 561 57 593 91
rect 631 57 663 91
rect 663 57 665 91
rect -1046 -48 -1012 -14
rect 1012 -48 1046 -14
<< metal1 >>
rect -701 91 701 97
rect -701 57 -665 91
rect -631 57 -593 91
rect -559 57 -521 91
rect -487 57 -449 91
rect -415 57 -377 91
rect -343 57 -305 91
rect -271 57 -233 91
rect -199 57 -161 91
rect -127 57 -89 91
rect -55 57 -17 91
rect 17 57 55 91
rect 89 57 127 91
rect 161 57 199 91
rect 233 57 271 91
rect 305 57 343 91
rect 377 57 415 91
rect 449 57 487 91
rect 521 57 559 91
rect 593 57 631 91
rect 665 57 701 91
rect -701 51 701 57
rect -1052 -14 -1006 8
rect -1052 -48 -1046 -14
rect -1012 -48 -1006 -14
rect -1052 -70 -1006 -48
rect 1006 -14 1052 8
rect 1006 -48 1012 -14
rect 1046 -48 1052 -14
rect 1006 -70 1052 -48
<< end >>
