magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -134 -107 134 45
<< nmoslvt >>
rect -50 -81 50 19
<< ndiff >>
rect -108 -14 -50 19
rect -108 -48 -96 -14
rect -62 -48 -50 -14
rect -108 -81 -50 -48
rect 50 -14 108 19
rect 50 -48 62 -14
rect 96 -48 108 -14
rect 50 -81 108 -48
<< ndiffc >>
rect -96 -48 -62 -14
rect 62 -48 96 -14
<< poly >>
rect -50 91 50 107
rect -50 57 -17 91
rect 17 57 50 91
rect -50 19 50 57
rect -50 -107 50 -81
<< polycont >>
rect -17 57 17 91
<< locali >>
rect -50 57 -17 91
rect 17 57 50 91
rect -96 -14 -62 23
rect -96 -85 -62 -48
rect 62 -14 96 23
rect 62 -85 96 -48
<< viali >>
rect -17 57 17 91
rect -96 -48 -62 -14
rect 62 -48 96 -14
<< metal1 >>
rect -46 91 46 97
rect -46 57 -17 91
rect 17 57 46 91
rect -46 51 46 57
rect -102 -14 -56 19
rect -102 -48 -96 -14
rect -62 -48 -56 -14
rect -102 -81 -56 -48
rect 56 -14 102 19
rect 56 -48 62 -14
rect 96 -48 102 -14
rect 56 -81 102 -48
<< end >>
