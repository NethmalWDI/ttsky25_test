magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -194 -198 194 164
<< pmoslvt >>
rect -100 -136 100 64
<< pdiff >>
rect -158 15 -100 64
rect -158 -19 -146 15
rect -112 -19 -100 15
rect -158 -53 -100 -19
rect -158 -87 -146 -53
rect -112 -87 -100 -53
rect -158 -136 -100 -87
rect 100 15 158 64
rect 100 -19 112 15
rect 146 -19 158 15
rect 100 -53 158 -19
rect 100 -87 112 -53
rect 146 -87 158 -53
rect 100 -136 158 -87
<< pdiffc >>
rect -146 -19 -112 15
rect -146 -87 -112 -53
rect 112 -19 146 15
rect 112 -87 146 -53
<< poly >>
rect -75 145 75 161
rect -75 128 -51 145
rect -100 111 -51 128
rect -17 111 17 145
rect 51 128 75 145
rect 51 111 100 128
rect -100 64 100 111
rect -100 -162 100 -136
<< polycont >>
rect -51 111 -17 145
rect 17 111 51 145
<< locali >>
rect -75 111 -53 145
rect -17 111 17 145
rect 53 111 75 145
rect -146 17 -112 42
rect -146 -53 -112 -19
rect -146 -114 -112 -89
rect 112 17 146 42
rect 112 -53 146 -19
rect 112 -114 146 -89
<< viali >>
rect -53 111 -51 145
rect -51 111 -19 145
rect 19 111 51 145
rect 51 111 53 145
rect -146 15 -112 17
rect -146 -17 -112 15
rect -146 -87 -112 -55
rect -146 -89 -112 -87
rect 112 15 146 17
rect 112 -17 146 15
rect 112 -87 146 -55
rect 112 -89 146 -87
<< metal1 >>
rect -71 145 71 151
rect -71 111 -53 145
rect -19 111 19 145
rect 53 111 71 145
rect -71 105 71 111
rect -152 17 -106 38
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -110 -106 -89
rect 106 17 152 38
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -110 152 -89
<< end >>
