magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< metal1 >>
rect 8900 7440 8980 7450
rect 8900 7436 9170 7440
rect 8900 7384 8914 7436
rect 8966 7426 9170 7436
rect 8966 7384 9114 7426
rect 8900 7380 9114 7384
rect 8900 7370 8980 7380
rect 9110 7374 9114 7380
rect 9166 7374 9170 7426
rect 9110 7360 9170 7374
<< via1 >>
rect 8914 7384 8966 7436
rect 9114 7374 9166 7426
<< metal2 >>
rect 9280 7530 9360 7540
rect 9010 7528 9360 7530
rect 9010 7472 9292 7528
rect 9348 7472 9360 7528
rect 9010 7470 9360 7472
rect 8900 7438 8980 7450
rect 8900 7382 8912 7438
rect 8968 7382 8980 7438
rect 8900 7370 8980 7382
rect 8796 4842 8876 4852
rect 9010 4842 9070 7470
rect 9280 7460 9360 7470
rect 9110 7426 9170 7440
rect 9110 7374 9114 7426
rect 9166 7374 9170 7426
rect 9110 5042 9170 7374
rect 9110 4982 9466 5042
rect 8796 4840 9070 4842
rect 8796 4784 8808 4840
rect 8864 4784 9070 4840
rect 8796 4782 9070 4784
rect 9406 4782 9466 4982
rect 8796 4772 8876 4782
rect 9406 4770 9486 4782
rect 9406 4714 9418 4770
rect 9474 4714 9486 4770
rect 9406 4702 9486 4714
<< via2 >>
rect 9292 7472 9348 7528
rect 8912 7436 8968 7438
rect 8912 7384 8914 7436
rect 8914 7384 8966 7436
rect 8966 7384 8968 7436
rect 8912 7382 8968 7384
rect 8808 4784 8864 4840
rect 9418 4714 9474 4770
<< metal3 >>
rect 14860 9248 14881 9252
rect 13920 7890 14940 7892
rect 13930 7602 14940 7890
rect 13930 7600 13960 7602
rect 9290 7528 9350 7530
rect 9290 7472 9292 7528
rect 9348 7472 9350 7528
rect 9290 7470 9350 7472
rect 8900 7438 8980 7450
rect 8900 7382 8912 7438
rect 8968 7382 8980 7438
rect 8900 7370 8980 7382
rect 13920 4962 14940 5270
rect 15230 5227 15320 5240
rect 15230 5163 15243 5227
rect 15307 5163 15320 5227
rect 15230 5150 15320 5163
rect 13920 4960 13960 4962
rect 8796 4840 8876 4852
rect 8796 4784 8808 4840
rect 8864 4784 8876 4840
rect 8796 4772 8876 4784
rect 9406 4770 9486 4782
rect 9406 4714 9418 4770
rect 9474 4714 9486 4770
rect 9406 4702 9486 4714
rect 15230 2500 15290 5150
rect 15230 2487 15320 2500
rect 15230 2423 15243 2487
rect 15307 2423 15320 2487
rect 15230 2410 15320 2423
<< via3 >>
rect 15243 5163 15307 5227
rect 15243 2423 15307 2487
<< metal4 >>
rect 1010 9250 13870 9252
rect 14040 9250 14881 9252
rect 1010 9248 14881 9250
rect 1010 8880 14861 9248
rect 1010 8772 1250 8880
rect 1010 7920 1252 8772
rect 1010 7610 1250 7920
rect 15070 7850 15510 7890
rect 8940 7830 15510 7850
rect 8940 7790 15130 7830
rect 15410 7790 15510 7830
rect 1010 5320 1252 7610
rect 4230 7608 4410 7610
rect 4230 7512 4670 7608
rect 4230 7510 4410 7512
rect 6650 7510 6970 7610
rect 8940 7520 9000 7790
rect 13560 7670 15130 7730
rect 11490 7608 11670 7610
rect 11290 7512 11670 7608
rect 13560 7520 13620 7670
rect 15070 7650 15130 7670
rect 15410 7650 15510 7690
rect 11490 7510 11670 7512
rect 14000 7210 14150 7610
rect 15070 7590 15510 7650
rect 4220 5320 4720 5430
rect 6550 5320 7050 5450
rect 8870 5352 8930 5360
rect 1010 4970 1250 5320
rect 8770 5094 8930 5352
rect 11230 5320 11710 5440
rect 13490 5229 13591 5319
rect 13490 5227 15450 5229
rect 13490 5163 15243 5227
rect 15307 5163 15450 5227
rect 13490 5160 15450 5163
rect 15230 5142 15450 5160
rect 8770 5032 15110 5094
rect 15050 5010 15110 5032
rect 15350 5010 15450 5032
rect 1010 1059 1252 4970
rect 4290 4870 4670 4970
rect 6650 4870 6970 4970
rect 11290 4870 11690 4970
rect 14000 4560 14170 4960
rect 15050 4950 15450 5010
rect 4210 2680 4710 2800
rect 6540 2680 7040 2800
rect 8770 2472 8930 2692
rect 11240 2680 11720 2780
rect 13490 2590 13550 2730
rect 15050 2590 15110 4950
rect 15350 4932 15450 4950
rect 13490 2530 15110 2590
rect 15230 2487 15320 2500
rect 8770 2470 8990 2472
rect 15230 2470 15243 2487
rect 8770 2423 15243 2470
rect 15307 2423 15320 2487
rect 8770 2412 15320 2423
rect 8930 2410 15320 2412
rect 2390 1980 2490 2290
rect 4700 1970 4800 2280
rect 7010 1970 7110 2280
rect 9320 1970 9420 2280
rect 11630 1970 11730 2280
rect 14000 1930 14160 2270
rect 2370 1160 2400 1162
rect 1870 1062 14860 1160
rect 1870 1060 2020 1062
rect 2350 1060 14860 1062
use sky130_fd_pr__cap_mim_m3_1_B9M9HY  sky130_fd_pr__cap_mim_m3_1_B9M9HY_0
timestamp 1757161594
transform 0 -1 3310 1 0 6426
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_0
timestamp 1757161594
transform 0 -1 3310 1 0 1666
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_1
timestamp 1757161594
transform 0 -1 5640 1 0 1666
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_2
timestamp 1757161594
transform 0 -1 7970 1 0 1666
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_3
timestamp 1757161594
transform 0 -1 10300 1 0 1666
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_4
timestamp 1757161594
transform 0 -1 12630 1 0 1666
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_5
timestamp 1757161594
transform 0 -1 12630 1 0 8566
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_6
timestamp 1757161594
transform 0 -1 10300 1 0 8566
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_7
timestamp 1757161594
transform 0 -1 7970 1 0 8566
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_8
timestamp 1757161594
transform 0 -1 5640 1 0 8566
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_DP2CMY  sky130_fd_pr__cap_mim_m3_1_DP2CMY_9
timestamp 1757161594
transform 0 -1 3310 1 0 8566
box -686 -1040 686 1040
use sky130_fd_pr__cap_mim_m3_1_G6WD7P  sky130_fd_pr__cap_mim_m3_1_G6WD7P_0
timestamp 1757161594
transform 0 -1 1440 1 0 1666
box -686 -540 686 540
use sky130_fd_pr__cap_mim_m3_1_G6WD7P  sky130_fd_pr__cap_mim_m3_1_G6WD7P_1
timestamp 1757161594
transform 0 -1 14460 1 0 1666
box -686 -540 686 540
use sky130_fd_pr__cap_mim_m3_1_G6WD7P  sky130_fd_pr__cap_mim_m3_1_G6WD7P_2
timestamp 1757161594
transform 0 -1 1440 1 0 8566
box -686 -540 686 540
use sky130_fd_pr__cap_mim_m3_1_G6WD7P  sky130_fd_pr__cap_mim_m3_1_G6WD7P_3
timestamp 1757161594
transform 0 -1 14460 1 0 8566
box -686 -540 686 540
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_1
timestamp 1757161594
transform 0 -1 10300 1 0 3786
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_3
timestamp 1757161594
transform 0 -1 5640 1 0 3786
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_4
timestamp 1757161594
transform 0 -1 7970 1 0 3786
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_5
timestamp 1757161594
transform 0 -1 3310 1 0 3786
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_6
timestamp 1757161594
transform 0 -1 12630 1 0 3786
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_15
timestamp 1757161594
transform 0 -1 5640 1 0 6426
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_17
timestamp 1757161594
transform 0 -1 7970 1 0 6426
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_18
timestamp 1757161594
transform 0 -1 12630 1 0 6426
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_GQMTM9  sky130_fd_pr__cap_mim_m3_1_GQMTM9_19
timestamp 1757161594
transform 0 -1 10300 1 0 6426
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_MYAC2F  sky130_fd_pr__cap_mim_m3_1_MYAC2F_0
timestamp 1757161594
transform 0 -1 14460 1 0 6426
box -1186 -540 1186 540
use sky130_fd_pr__cap_mim_m3_1_MYAC2F  sky130_fd_pr__cap_mim_m3_1_MYAC2F_1
timestamp 1757161594
transform 0 -1 14460 1 0 3786
box -1186 -540 1186 540
use sky130_fd_pr__cap_mim_m3_1_MYAC2F  sky130_fd_pr__cap_mim_m3_1_MYAC2F_2
timestamp 1757161594
transform 0 -1 1440 1 0 3786
box -1186 -540 1186 540
use sky130_fd_pr__cap_mim_m3_1_MYAC2F  sky130_fd_pr__cap_mim_m3_1_MYAC2F_3
timestamp 1757161594
transform 0 -1 1440 1 0 6426
box -1186 -540 1186 540
<< end >>
