magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< error_s >>
rect 6467 5290 6577 5358
rect 6707 5290 6817 5358
rect 6467 5190 6635 5290
rect 6707 5190 6875 5290
rect 6193 -573 6893 -336
rect 6447 -590 6557 -573
rect 6697 -590 6807 -573
rect 6557 -690 6615 -590
rect 6697 -690 6865 -590
<< nwell >>
rect 6467 5190 6577 5290
rect 6707 5190 6817 5290
rect 57 5163 237 5170
rect -313 -573 6893 5163
rect 6447 -690 6557 -590
rect 6697 -690 6807 -590
<< nsubdiff >>
rect -277 5093 -195 5127
rect -161 5093 -127 5127
rect -93 5093 -59 5127
rect -25 5093 9 5127
rect 43 5093 77 5127
rect 111 5093 145 5127
rect 179 5093 213 5127
rect 247 5093 281 5127
rect 315 5093 349 5127
rect 383 5093 417 5127
rect 451 5093 485 5127
rect 519 5093 553 5127
rect 587 5093 621 5127
rect 655 5093 689 5127
rect 723 5093 757 5127
rect 791 5093 825 5127
rect 859 5093 893 5127
rect 927 5093 961 5127
rect 995 5093 1029 5127
rect 1063 5093 1097 5127
rect 1131 5093 1165 5127
rect 1199 5093 1233 5127
rect 1267 5093 1301 5127
rect 1335 5093 1369 5127
rect 1403 5093 1437 5127
rect 1471 5093 1505 5127
rect 1539 5093 1573 5127
rect 1607 5093 1641 5127
rect 1675 5093 1709 5127
rect 1743 5093 1777 5127
rect 1811 5093 1845 5127
rect 1879 5093 1913 5127
rect 1947 5093 1981 5127
rect 2015 5093 2049 5127
rect 2083 5093 2117 5127
rect 2151 5093 2185 5127
rect 2219 5093 2253 5127
rect 2287 5093 2321 5127
rect 2355 5093 2389 5127
rect 2423 5093 2457 5127
rect 2491 5093 2525 5127
rect 2559 5093 2593 5127
rect 2627 5093 2661 5127
rect 2695 5093 2729 5127
rect 2763 5093 2797 5127
rect 2831 5093 2865 5127
rect 2899 5093 2933 5127
rect 2967 5093 3001 5127
rect 3035 5093 3069 5127
rect 3103 5093 3137 5127
rect 3171 5093 3205 5127
rect 3239 5093 3273 5127
rect 3307 5093 3341 5127
rect 3375 5093 3409 5127
rect 3443 5093 3477 5127
rect 3511 5093 3545 5127
rect 3579 5093 3613 5127
rect 3647 5093 3681 5127
rect 3715 5093 3749 5127
rect 3783 5093 3817 5127
rect 3851 5093 3885 5127
rect 3919 5093 3953 5127
rect 3987 5093 4021 5127
rect 4055 5093 4089 5127
rect 4123 5093 4157 5127
rect 4191 5093 4225 5127
rect 4259 5093 4293 5127
rect 4327 5093 4361 5127
rect 4395 5093 4429 5127
rect 4463 5093 4497 5127
rect 4531 5093 4565 5127
rect 4599 5093 4633 5127
rect 4667 5093 4701 5127
rect 4735 5093 4769 5127
rect 4803 5093 4837 5127
rect 4871 5093 4905 5127
rect 4939 5093 4973 5127
rect 5007 5093 5041 5127
rect 5075 5093 5109 5127
rect 5143 5093 5177 5127
rect 5211 5093 5245 5127
rect 5279 5093 5313 5127
rect 5347 5093 5381 5127
rect 5415 5093 5449 5127
rect 5483 5093 5517 5127
rect 5551 5093 5585 5127
rect 5619 5093 5653 5127
rect 5687 5093 5721 5127
rect 5755 5093 5789 5127
rect 5823 5093 5857 5127
rect 5891 5093 5925 5127
rect 5959 5093 5993 5127
rect 6027 5093 6061 5127
rect 6095 5093 6129 5127
rect 6163 5093 6197 5127
rect 6231 5093 6265 5127
rect 6299 5093 6333 5127
rect 6367 5093 6401 5127
rect 6435 5093 6469 5127
rect 6503 5093 6537 5127
rect 6571 5093 6605 5127
rect 6639 5093 6673 5127
rect 6707 5093 6741 5127
rect 6775 5093 6857 5127
rect -277 5066 -243 5093
rect -277 4998 -243 5032
rect -277 4930 -243 4964
rect -277 4862 -243 4896
rect -277 4794 -243 4828
rect -277 4726 -243 4760
rect -277 4658 -243 4692
rect -277 4590 -243 4624
rect -277 4522 -243 4556
rect -277 4454 -243 4488
rect -277 4386 -243 4420
rect -277 4318 -243 4352
rect -277 4250 -243 4284
rect -277 4182 -243 4216
rect -277 4114 -243 4148
rect -277 4046 -243 4080
rect -277 3978 -243 4012
rect -277 3910 -243 3944
rect -277 3842 -243 3876
rect -277 3774 -243 3808
rect -277 3706 -243 3740
rect -277 3638 -243 3672
rect -277 3570 -243 3604
rect -277 3502 -243 3536
rect -277 3434 -243 3468
rect -277 3366 -243 3400
rect -277 3298 -243 3332
rect -277 3230 -243 3264
rect -277 3162 -243 3196
rect -277 3094 -243 3128
rect -277 3026 -243 3060
rect -277 2958 -243 2992
rect -277 2890 -243 2924
rect -277 2822 -243 2856
rect -277 2754 -243 2788
rect -277 2686 -243 2720
rect -277 2618 -243 2652
rect -277 2550 -243 2584
rect -277 2482 -243 2516
rect -277 2414 -243 2448
rect -277 2346 -243 2380
rect -277 2278 -243 2312
rect -277 2210 -243 2244
rect -277 2142 -243 2176
rect -277 2074 -243 2108
rect -277 2006 -243 2040
rect -277 1938 -243 1972
rect -277 1870 -243 1904
rect -277 1802 -243 1836
rect -277 1734 -243 1768
rect -277 1666 -243 1700
rect -277 1598 -243 1632
rect -277 1530 -243 1564
rect -277 1462 -243 1496
rect -277 1394 -243 1428
rect -277 1326 -243 1360
rect -277 1258 -243 1292
rect -277 1190 -243 1224
rect -277 1122 -243 1156
rect -277 1054 -243 1088
rect -277 986 -243 1020
rect -277 918 -243 952
rect -277 850 -243 884
rect -277 782 -243 816
rect -277 714 -243 748
rect -277 646 -243 680
rect -277 578 -243 612
rect -277 510 -243 544
rect -277 442 -243 476
rect -277 374 -243 408
rect -277 306 -243 340
rect -277 238 -243 272
rect -277 170 -243 204
rect -277 102 -243 136
rect -277 34 -243 68
rect -277 -34 -243 0
rect -277 -102 -243 -68
rect -277 -170 -243 -136
rect -277 -238 -243 -204
rect -277 -306 -243 -272
rect -277 -374 -243 -340
rect -277 -442 -243 -408
rect -277 -503 -243 -476
rect 6823 5066 6857 5093
rect 6823 4998 6857 5032
rect 6823 4930 6857 4964
rect 6823 4862 6857 4896
rect 6823 4794 6857 4828
rect 6823 4726 6857 4760
rect 6823 4658 6857 4692
rect 6823 4590 6857 4624
rect 6823 4522 6857 4556
rect 6823 4454 6857 4488
rect 6823 4386 6857 4420
rect 6823 4318 6857 4352
rect 6823 4250 6857 4284
rect 6823 4182 6857 4216
rect 6823 4114 6857 4148
rect 6823 4046 6857 4080
rect 6823 3978 6857 4012
rect 6823 3910 6857 3944
rect 6823 3842 6857 3876
rect 6823 3774 6857 3808
rect 6823 3706 6857 3740
rect 6823 3638 6857 3672
rect 6823 3570 6857 3604
rect 6823 3502 6857 3536
rect 6823 3434 6857 3468
rect 6823 3366 6857 3400
rect 6823 3298 6857 3332
rect 6823 3230 6857 3264
rect 6823 3162 6857 3196
rect 6823 3094 6857 3128
rect 6823 3026 6857 3060
rect 6823 2958 6857 2992
rect 6823 2890 6857 2924
rect 6823 2822 6857 2856
rect 6823 2754 6857 2788
rect 6823 2686 6857 2720
rect 6823 2618 6857 2652
rect 6823 2550 6857 2584
rect 6823 2482 6857 2516
rect 6823 2414 6857 2448
rect 6823 2346 6857 2380
rect 6823 2278 6857 2312
rect 6823 2210 6857 2244
rect 6823 2142 6857 2176
rect 6823 2074 6857 2108
rect 6823 2006 6857 2040
rect 6823 1938 6857 1972
rect 6823 1870 6857 1904
rect 6823 1802 6857 1836
rect 6823 1734 6857 1768
rect 6823 1666 6857 1700
rect 6823 1598 6857 1632
rect 6823 1530 6857 1564
rect 6823 1462 6857 1496
rect 6823 1394 6857 1428
rect 6823 1326 6857 1360
rect 6823 1258 6857 1292
rect 6823 1190 6857 1224
rect 6823 1122 6857 1156
rect 6823 1054 6857 1088
rect 6823 986 6857 1020
rect 6823 918 6857 952
rect 6823 850 6857 884
rect 6823 782 6857 816
rect 6823 714 6857 748
rect 6823 646 6857 680
rect 6823 578 6857 612
rect 6823 510 6857 544
rect 6823 442 6857 476
rect 6823 374 6857 408
rect 6823 306 6857 340
rect 6823 238 6857 272
rect 6823 170 6857 204
rect 6823 102 6857 136
rect 6823 34 6857 68
rect 6823 -34 6857 0
rect 6823 -102 6857 -68
rect 6823 -170 6857 -136
rect 6823 -238 6857 -204
rect 6823 -306 6857 -272
rect 6823 -374 6857 -340
rect 6823 -442 6857 -408
rect 6823 -503 6857 -476
rect -277 -537 -195 -503
rect -161 -537 -127 -503
rect -93 -537 -59 -503
rect -25 -537 9 -503
rect 43 -537 77 -503
rect 111 -537 145 -503
rect 179 -537 213 -503
rect 247 -537 281 -503
rect 315 -537 349 -503
rect 383 -537 417 -503
rect 451 -537 485 -503
rect 519 -537 553 -503
rect 587 -537 621 -503
rect 655 -537 689 -503
rect 723 -537 757 -503
rect 791 -537 825 -503
rect 859 -537 893 -503
rect 927 -537 961 -503
rect 995 -537 1029 -503
rect 1063 -537 1097 -503
rect 1131 -537 1165 -503
rect 1199 -537 1233 -503
rect 1267 -537 1301 -503
rect 1335 -537 1369 -503
rect 1403 -537 1437 -503
rect 1471 -537 1505 -503
rect 1539 -537 1573 -503
rect 1607 -537 1641 -503
rect 1675 -537 1709 -503
rect 1743 -537 1777 -503
rect 1811 -537 1845 -503
rect 1879 -537 1913 -503
rect 1947 -537 1981 -503
rect 2015 -537 2049 -503
rect 2083 -537 2117 -503
rect 2151 -537 2185 -503
rect 2219 -537 2253 -503
rect 2287 -537 2321 -503
rect 2355 -537 2389 -503
rect 2423 -537 2457 -503
rect 2491 -537 2525 -503
rect 2559 -537 2593 -503
rect 2627 -537 2661 -503
rect 2695 -537 2729 -503
rect 2763 -537 2797 -503
rect 2831 -537 2865 -503
rect 2899 -537 2933 -503
rect 2967 -537 3001 -503
rect 3035 -537 3069 -503
rect 3103 -537 3137 -503
rect 3171 -537 3205 -503
rect 3239 -537 3273 -503
rect 3307 -537 3341 -503
rect 3375 -537 3409 -503
rect 3443 -537 3477 -503
rect 3511 -537 3545 -503
rect 3579 -537 3613 -503
rect 3647 -537 3681 -503
rect 3715 -537 3749 -503
rect 3783 -537 3817 -503
rect 3851 -537 3885 -503
rect 3919 -537 3953 -503
rect 3987 -537 4021 -503
rect 4055 -537 4089 -503
rect 4123 -537 4157 -503
rect 4191 -537 4225 -503
rect 4259 -537 4293 -503
rect 4327 -537 4361 -503
rect 4395 -537 4429 -503
rect 4463 -537 4497 -503
rect 4531 -537 4565 -503
rect 4599 -537 4633 -503
rect 4667 -537 4701 -503
rect 4735 -537 4769 -503
rect 4803 -537 4837 -503
rect 4871 -537 4905 -503
rect 4939 -537 4973 -503
rect 5007 -537 5041 -503
rect 5075 -537 5109 -503
rect 5143 -537 5177 -503
rect 5211 -537 5245 -503
rect 5279 -537 5313 -503
rect 5347 -537 5381 -503
rect 5415 -537 5449 -503
rect 5483 -537 5517 -503
rect 5551 -537 5585 -503
rect 5619 -537 5653 -503
rect 5687 -537 5721 -503
rect 5755 -537 5789 -503
rect 5823 -537 5857 -503
rect 5891 -537 5925 -503
rect 5959 -537 5993 -503
rect 6027 -537 6061 -503
rect 6095 -537 6129 -503
rect 6163 -537 6197 -503
rect 6231 -537 6265 -503
rect 6299 -537 6333 -503
rect 6367 -537 6401 -503
rect 6435 -537 6469 -503
rect 6503 -537 6537 -503
rect 6571 -537 6605 -503
rect 6639 -537 6673 -503
rect 6707 -537 6741 -503
rect 6775 -537 6857 -503
<< nsubdiffcont >>
rect -195 5093 -161 5127
rect -127 5093 -93 5127
rect -59 5093 -25 5127
rect 9 5093 43 5127
rect 77 5093 111 5127
rect 145 5093 179 5127
rect 213 5093 247 5127
rect 281 5093 315 5127
rect 349 5093 383 5127
rect 417 5093 451 5127
rect 485 5093 519 5127
rect 553 5093 587 5127
rect 621 5093 655 5127
rect 689 5093 723 5127
rect 757 5093 791 5127
rect 825 5093 859 5127
rect 893 5093 927 5127
rect 961 5093 995 5127
rect 1029 5093 1063 5127
rect 1097 5093 1131 5127
rect 1165 5093 1199 5127
rect 1233 5093 1267 5127
rect 1301 5093 1335 5127
rect 1369 5093 1403 5127
rect 1437 5093 1471 5127
rect 1505 5093 1539 5127
rect 1573 5093 1607 5127
rect 1641 5093 1675 5127
rect 1709 5093 1743 5127
rect 1777 5093 1811 5127
rect 1845 5093 1879 5127
rect 1913 5093 1947 5127
rect 1981 5093 2015 5127
rect 2049 5093 2083 5127
rect 2117 5093 2151 5127
rect 2185 5093 2219 5127
rect 2253 5093 2287 5127
rect 2321 5093 2355 5127
rect 2389 5093 2423 5127
rect 2457 5093 2491 5127
rect 2525 5093 2559 5127
rect 2593 5093 2627 5127
rect 2661 5093 2695 5127
rect 2729 5093 2763 5127
rect 2797 5093 2831 5127
rect 2865 5093 2899 5127
rect 2933 5093 2967 5127
rect 3001 5093 3035 5127
rect 3069 5093 3103 5127
rect 3137 5093 3171 5127
rect 3205 5093 3239 5127
rect 3273 5093 3307 5127
rect 3341 5093 3375 5127
rect 3409 5093 3443 5127
rect 3477 5093 3511 5127
rect 3545 5093 3579 5127
rect 3613 5093 3647 5127
rect 3681 5093 3715 5127
rect 3749 5093 3783 5127
rect 3817 5093 3851 5127
rect 3885 5093 3919 5127
rect 3953 5093 3987 5127
rect 4021 5093 4055 5127
rect 4089 5093 4123 5127
rect 4157 5093 4191 5127
rect 4225 5093 4259 5127
rect 4293 5093 4327 5127
rect 4361 5093 4395 5127
rect 4429 5093 4463 5127
rect 4497 5093 4531 5127
rect 4565 5093 4599 5127
rect 4633 5093 4667 5127
rect 4701 5093 4735 5127
rect 4769 5093 4803 5127
rect 4837 5093 4871 5127
rect 4905 5093 4939 5127
rect 4973 5093 5007 5127
rect 5041 5093 5075 5127
rect 5109 5093 5143 5127
rect 5177 5093 5211 5127
rect 5245 5093 5279 5127
rect 5313 5093 5347 5127
rect 5381 5093 5415 5127
rect 5449 5093 5483 5127
rect 5517 5093 5551 5127
rect 5585 5093 5619 5127
rect 5653 5093 5687 5127
rect 5721 5093 5755 5127
rect 5789 5093 5823 5127
rect 5857 5093 5891 5127
rect 5925 5093 5959 5127
rect 5993 5093 6027 5127
rect 6061 5093 6095 5127
rect 6129 5093 6163 5127
rect 6197 5093 6231 5127
rect 6265 5093 6299 5127
rect 6333 5093 6367 5127
rect 6401 5093 6435 5127
rect 6469 5093 6503 5127
rect 6537 5093 6571 5127
rect 6605 5093 6639 5127
rect 6673 5093 6707 5127
rect 6741 5093 6775 5127
rect -277 5032 -243 5066
rect -277 4964 -243 4998
rect -277 4896 -243 4930
rect -277 4828 -243 4862
rect -277 4760 -243 4794
rect -277 4692 -243 4726
rect -277 4624 -243 4658
rect -277 4556 -243 4590
rect -277 4488 -243 4522
rect -277 4420 -243 4454
rect -277 4352 -243 4386
rect -277 4284 -243 4318
rect -277 4216 -243 4250
rect -277 4148 -243 4182
rect -277 4080 -243 4114
rect -277 4012 -243 4046
rect -277 3944 -243 3978
rect -277 3876 -243 3910
rect -277 3808 -243 3842
rect -277 3740 -243 3774
rect -277 3672 -243 3706
rect -277 3604 -243 3638
rect -277 3536 -243 3570
rect -277 3468 -243 3502
rect -277 3400 -243 3434
rect -277 3332 -243 3366
rect -277 3264 -243 3298
rect -277 3196 -243 3230
rect -277 3128 -243 3162
rect -277 3060 -243 3094
rect -277 2992 -243 3026
rect -277 2924 -243 2958
rect -277 2856 -243 2890
rect -277 2788 -243 2822
rect -277 2720 -243 2754
rect -277 2652 -243 2686
rect -277 2584 -243 2618
rect -277 2516 -243 2550
rect -277 2448 -243 2482
rect -277 2380 -243 2414
rect -277 2312 -243 2346
rect -277 2244 -243 2278
rect -277 2176 -243 2210
rect -277 2108 -243 2142
rect -277 2040 -243 2074
rect -277 1972 -243 2006
rect -277 1904 -243 1938
rect -277 1836 -243 1870
rect -277 1768 -243 1802
rect -277 1700 -243 1734
rect -277 1632 -243 1666
rect -277 1564 -243 1598
rect -277 1496 -243 1530
rect -277 1428 -243 1462
rect -277 1360 -243 1394
rect -277 1292 -243 1326
rect -277 1224 -243 1258
rect -277 1156 -243 1190
rect -277 1088 -243 1122
rect -277 1020 -243 1054
rect -277 952 -243 986
rect -277 884 -243 918
rect -277 816 -243 850
rect -277 748 -243 782
rect -277 680 -243 714
rect -277 612 -243 646
rect -277 544 -243 578
rect -277 476 -243 510
rect -277 408 -243 442
rect -277 340 -243 374
rect -277 272 -243 306
rect -277 204 -243 238
rect -277 136 -243 170
rect -277 68 -243 102
rect -277 0 -243 34
rect -277 -68 -243 -34
rect -277 -136 -243 -102
rect -277 -204 -243 -170
rect -277 -272 -243 -238
rect -277 -340 -243 -306
rect -277 -408 -243 -374
rect -277 -476 -243 -442
rect 6823 5032 6857 5066
rect 6823 4964 6857 4998
rect 6823 4896 6857 4930
rect 6823 4828 6857 4862
rect 6823 4760 6857 4794
rect 6823 4692 6857 4726
rect 6823 4624 6857 4658
rect 6823 4556 6857 4590
rect 6823 4488 6857 4522
rect 6823 4420 6857 4454
rect 6823 4352 6857 4386
rect 6823 4284 6857 4318
rect 6823 4216 6857 4250
rect 6823 4148 6857 4182
rect 6823 4080 6857 4114
rect 6823 4012 6857 4046
rect 6823 3944 6857 3978
rect 6823 3876 6857 3910
rect 6823 3808 6857 3842
rect 6823 3740 6857 3774
rect 6823 3672 6857 3706
rect 6823 3604 6857 3638
rect 6823 3536 6857 3570
rect 6823 3468 6857 3502
rect 6823 3400 6857 3434
rect 6823 3332 6857 3366
rect 6823 3264 6857 3298
rect 6823 3196 6857 3230
rect 6823 3128 6857 3162
rect 6823 3060 6857 3094
rect 6823 2992 6857 3026
rect 6823 2924 6857 2958
rect 6823 2856 6857 2890
rect 6823 2788 6857 2822
rect 6823 2720 6857 2754
rect 6823 2652 6857 2686
rect 6823 2584 6857 2618
rect 6823 2516 6857 2550
rect 6823 2448 6857 2482
rect 6823 2380 6857 2414
rect 6823 2312 6857 2346
rect 6823 2244 6857 2278
rect 6823 2176 6857 2210
rect 6823 2108 6857 2142
rect 6823 2040 6857 2074
rect 6823 1972 6857 2006
rect 6823 1904 6857 1938
rect 6823 1836 6857 1870
rect 6823 1768 6857 1802
rect 6823 1700 6857 1734
rect 6823 1632 6857 1666
rect 6823 1564 6857 1598
rect 6823 1496 6857 1530
rect 6823 1428 6857 1462
rect 6823 1360 6857 1394
rect 6823 1292 6857 1326
rect 6823 1224 6857 1258
rect 6823 1156 6857 1190
rect 6823 1088 6857 1122
rect 6823 1020 6857 1054
rect 6823 952 6857 986
rect 6823 884 6857 918
rect 6823 816 6857 850
rect 6823 748 6857 782
rect 6823 680 6857 714
rect 6823 612 6857 646
rect 6823 544 6857 578
rect 6823 476 6857 510
rect 6823 408 6857 442
rect 6823 340 6857 374
rect 6823 272 6857 306
rect 6823 204 6857 238
rect 6823 136 6857 170
rect 6823 68 6857 102
rect 6823 0 6857 34
rect 6823 -68 6857 -34
rect 6823 -136 6857 -102
rect 6823 -204 6857 -170
rect 6823 -272 6857 -238
rect 6823 -340 6857 -306
rect 6823 -408 6857 -374
rect 6823 -476 6857 -442
rect -195 -537 -161 -503
rect -127 -537 -93 -503
rect -59 -537 -25 -503
rect 9 -537 43 -503
rect 77 -537 111 -503
rect 145 -537 179 -503
rect 213 -537 247 -503
rect 281 -537 315 -503
rect 349 -537 383 -503
rect 417 -537 451 -503
rect 485 -537 519 -503
rect 553 -537 587 -503
rect 621 -537 655 -503
rect 689 -537 723 -503
rect 757 -537 791 -503
rect 825 -537 859 -503
rect 893 -537 927 -503
rect 961 -537 995 -503
rect 1029 -537 1063 -503
rect 1097 -537 1131 -503
rect 1165 -537 1199 -503
rect 1233 -537 1267 -503
rect 1301 -537 1335 -503
rect 1369 -537 1403 -503
rect 1437 -537 1471 -503
rect 1505 -537 1539 -503
rect 1573 -537 1607 -503
rect 1641 -537 1675 -503
rect 1709 -537 1743 -503
rect 1777 -537 1811 -503
rect 1845 -537 1879 -503
rect 1913 -537 1947 -503
rect 1981 -537 2015 -503
rect 2049 -537 2083 -503
rect 2117 -537 2151 -503
rect 2185 -537 2219 -503
rect 2253 -537 2287 -503
rect 2321 -537 2355 -503
rect 2389 -537 2423 -503
rect 2457 -537 2491 -503
rect 2525 -537 2559 -503
rect 2593 -537 2627 -503
rect 2661 -537 2695 -503
rect 2729 -537 2763 -503
rect 2797 -537 2831 -503
rect 2865 -537 2899 -503
rect 2933 -537 2967 -503
rect 3001 -537 3035 -503
rect 3069 -537 3103 -503
rect 3137 -537 3171 -503
rect 3205 -537 3239 -503
rect 3273 -537 3307 -503
rect 3341 -537 3375 -503
rect 3409 -537 3443 -503
rect 3477 -537 3511 -503
rect 3545 -537 3579 -503
rect 3613 -537 3647 -503
rect 3681 -537 3715 -503
rect 3749 -537 3783 -503
rect 3817 -537 3851 -503
rect 3885 -537 3919 -503
rect 3953 -537 3987 -503
rect 4021 -537 4055 -503
rect 4089 -537 4123 -503
rect 4157 -537 4191 -503
rect 4225 -537 4259 -503
rect 4293 -537 4327 -503
rect 4361 -537 4395 -503
rect 4429 -537 4463 -503
rect 4497 -537 4531 -503
rect 4565 -537 4599 -503
rect 4633 -537 4667 -503
rect 4701 -537 4735 -503
rect 4769 -537 4803 -503
rect 4837 -537 4871 -503
rect 4905 -537 4939 -503
rect 4973 -537 5007 -503
rect 5041 -537 5075 -503
rect 5109 -537 5143 -503
rect 5177 -537 5211 -503
rect 5245 -537 5279 -503
rect 5313 -537 5347 -503
rect 5381 -537 5415 -503
rect 5449 -537 5483 -503
rect 5517 -537 5551 -503
rect 5585 -537 5619 -503
rect 5653 -537 5687 -503
rect 5721 -537 5755 -503
rect 5789 -537 5823 -503
rect 5857 -537 5891 -503
rect 5925 -537 5959 -503
rect 5993 -537 6027 -503
rect 6061 -537 6095 -503
rect 6129 -537 6163 -503
rect 6197 -537 6231 -503
rect 6265 -537 6299 -503
rect 6333 -537 6367 -503
rect 6401 -537 6435 -503
rect 6469 -537 6503 -503
rect 6537 -537 6571 -503
rect 6605 -537 6639 -503
rect 6673 -537 6707 -503
rect 6741 -537 6775 -503
<< locali >>
rect -277 5093 -195 5127
rect -161 5093 -127 5127
rect -93 5093 -59 5127
rect -25 5093 9 5127
rect 43 5093 77 5127
rect 111 5093 145 5127
rect 179 5093 213 5127
rect 247 5093 281 5127
rect 315 5093 349 5127
rect 383 5093 417 5127
rect 451 5093 485 5127
rect 519 5093 553 5127
rect 587 5093 621 5127
rect 655 5093 689 5127
rect 723 5093 757 5127
rect 791 5093 825 5127
rect 859 5093 893 5127
rect 927 5093 961 5127
rect 995 5093 1029 5127
rect 1063 5093 1097 5127
rect 1131 5093 1165 5127
rect 1199 5093 1233 5127
rect 1267 5093 1301 5127
rect 1335 5093 1369 5127
rect 1403 5093 1437 5127
rect 1471 5093 1505 5127
rect 1539 5093 1573 5127
rect 1607 5093 1641 5127
rect 1675 5093 1709 5127
rect 1743 5093 1777 5127
rect 1811 5093 1845 5127
rect 1879 5093 1913 5127
rect 1947 5093 1981 5127
rect 2015 5093 2049 5127
rect 2083 5093 2117 5127
rect 2151 5093 2185 5127
rect 2219 5093 2253 5127
rect 2287 5093 2321 5127
rect 2355 5093 2389 5127
rect 2423 5093 2457 5127
rect 2491 5093 2525 5127
rect 2559 5093 2593 5127
rect 2627 5093 2661 5127
rect 2695 5093 2729 5127
rect 2763 5093 2797 5127
rect 2831 5093 2865 5127
rect 2899 5093 2933 5127
rect 2967 5093 3001 5127
rect 3035 5093 3069 5127
rect 3103 5093 3137 5127
rect 3171 5093 3205 5127
rect 3239 5093 3273 5127
rect 3307 5093 3341 5127
rect 3375 5093 3409 5127
rect 3443 5093 3477 5127
rect 3511 5093 3545 5127
rect 3579 5093 3613 5127
rect 3647 5093 3681 5127
rect 3715 5093 3749 5127
rect 3783 5093 3817 5127
rect 3851 5093 3885 5127
rect 3919 5093 3953 5127
rect 3987 5093 4021 5127
rect 4055 5093 4089 5127
rect 4123 5093 4157 5127
rect 4191 5093 4225 5127
rect 4259 5093 4293 5127
rect 4327 5093 4361 5127
rect 4395 5093 4429 5127
rect 4463 5093 4497 5127
rect 4531 5093 4565 5127
rect 4599 5093 4633 5127
rect 4667 5093 4701 5127
rect 4735 5093 4769 5127
rect 4803 5093 4837 5127
rect 4871 5093 4905 5127
rect 4939 5093 4973 5127
rect 5007 5093 5041 5127
rect 5075 5093 5109 5127
rect 5143 5093 5177 5127
rect 5211 5093 5245 5127
rect 5279 5093 5313 5127
rect 5347 5093 5381 5127
rect 5415 5093 5449 5127
rect 5483 5093 5517 5127
rect 5551 5093 5585 5127
rect 5619 5093 5653 5127
rect 5687 5093 5721 5127
rect 5755 5093 5789 5127
rect 5823 5093 5857 5127
rect 5891 5093 5925 5127
rect 5959 5093 5993 5127
rect 6027 5093 6061 5127
rect 6095 5093 6129 5127
rect 6163 5093 6197 5127
rect 6231 5093 6265 5127
rect 6299 5093 6333 5127
rect 6367 5093 6401 5127
rect 6435 5093 6469 5127
rect 6503 5093 6537 5127
rect 6571 5093 6605 5127
rect 6639 5093 6673 5127
rect 6707 5093 6741 5127
rect 6775 5093 6857 5127
rect -277 5066 -243 5093
rect -277 4998 -243 5032
rect -277 4930 -243 4964
rect -277 4862 -243 4896
rect -277 4794 -243 4828
rect -277 4726 -243 4760
rect -277 4658 -243 4692
rect -277 4590 -243 4624
rect -277 4522 -243 4556
rect -277 4454 -243 4488
rect -277 4386 -243 4420
rect -277 4318 -243 4352
rect -277 4250 -243 4284
rect -277 4182 -243 4216
rect -277 4114 -243 4148
rect -277 4046 -243 4080
rect -277 3978 -243 4012
rect -277 3910 -243 3944
rect -277 3842 -243 3876
rect -277 3774 -243 3808
rect -277 3706 -243 3740
rect -277 3638 -243 3672
rect -277 3570 -243 3604
rect -277 3502 -243 3536
rect -277 3434 -243 3468
rect -277 3366 -243 3400
rect -277 3298 -243 3332
rect -277 3230 -243 3264
rect -277 3162 -243 3196
rect -277 3094 -243 3128
rect -277 3026 -243 3060
rect -277 2958 -243 2992
rect -277 2890 -243 2924
rect -277 2822 -243 2856
rect -277 2754 -243 2788
rect -277 2686 -243 2720
rect -277 2618 -243 2652
rect -277 2550 -243 2584
rect -277 2482 -243 2516
rect -277 2414 -243 2448
rect -277 2346 -243 2380
rect -277 2278 -243 2312
rect -277 2210 -243 2244
rect -277 2142 -243 2176
rect -277 2074 -243 2108
rect -277 2006 -243 2040
rect -277 1938 -243 1972
rect -277 1870 -243 1904
rect -277 1802 -243 1836
rect -277 1734 -243 1768
rect -277 1666 -243 1700
rect -277 1598 -243 1632
rect -277 1530 -243 1564
rect -277 1462 -243 1496
rect -277 1394 -243 1428
rect -277 1326 -243 1360
rect -277 1258 -243 1292
rect -277 1190 -243 1224
rect -277 1122 -243 1156
rect -277 1054 -243 1088
rect -277 986 -243 1020
rect -277 918 -243 952
rect -277 850 -243 884
rect -277 782 -243 816
rect -277 714 -243 748
rect -277 646 -243 680
rect -277 578 -243 612
rect -277 510 -243 544
rect -277 442 -243 476
rect -277 374 -243 408
rect -277 306 -243 340
rect -277 238 -243 272
rect -277 170 -243 204
rect -277 102 -243 136
rect -277 34 -243 68
rect -277 -34 -243 0
rect -277 -102 -243 -68
rect -277 -170 -243 -136
rect -277 -238 -243 -204
rect -277 -306 -243 -272
rect -277 -374 -243 -340
rect -277 -442 -243 -408
rect -277 -503 -243 -476
rect 6823 5066 6857 5093
rect 6823 4998 6857 5032
rect 6823 4930 6857 4964
rect 6823 4862 6857 4896
rect 6823 4794 6857 4828
rect 6823 4726 6857 4760
rect 6823 4658 6857 4692
rect 6823 4590 6857 4624
rect 6823 4522 6857 4556
rect 6823 4454 6857 4488
rect 6823 4386 6857 4420
rect 6823 4318 6857 4352
rect 6823 4250 6857 4284
rect 6823 4182 6857 4216
rect 6823 4114 6857 4148
rect 6823 4046 6857 4080
rect 6823 3978 6857 4012
rect 6823 3910 6857 3944
rect 6823 3842 6857 3876
rect 6823 3774 6857 3808
rect 6823 3706 6857 3740
rect 6823 3638 6857 3672
rect 6823 3570 6857 3604
rect 6823 3502 6857 3536
rect 6823 3434 6857 3468
rect 6823 3366 6857 3400
rect 6823 3298 6857 3332
rect 6823 3230 6857 3264
rect 6823 3162 6857 3196
rect 6823 3094 6857 3128
rect 6823 3026 6857 3060
rect 6823 2958 6857 2992
rect 6823 2890 6857 2924
rect 6823 2822 6857 2856
rect 6823 2754 6857 2788
rect 6823 2686 6857 2720
rect 6823 2618 6857 2652
rect 6823 2550 6857 2584
rect 6823 2482 6857 2516
rect 6823 2414 6857 2448
rect 6823 2346 6857 2380
rect 6823 2278 6857 2312
rect 6823 2210 6857 2244
rect 6823 2142 6857 2176
rect 6823 2074 6857 2108
rect 6823 2006 6857 2040
rect 6823 1938 6857 1972
rect 6823 1870 6857 1904
rect 6823 1802 6857 1836
rect 6823 1734 6857 1768
rect 6823 1666 6857 1700
rect 6823 1598 6857 1632
rect 6823 1530 6857 1564
rect 6823 1462 6857 1496
rect 6823 1394 6857 1428
rect 6823 1326 6857 1360
rect 6823 1258 6857 1292
rect 6823 1190 6857 1224
rect 6823 1122 6857 1156
rect 6823 1054 6857 1088
rect 6823 986 6857 1020
rect 6823 918 6857 952
rect 6823 850 6857 884
rect 6823 782 6857 816
rect 6823 714 6857 748
rect 6823 646 6857 680
rect 6823 578 6857 612
rect 6823 510 6857 544
rect 6823 442 6857 476
rect 6823 374 6857 408
rect 6823 306 6857 340
rect 6823 238 6857 272
rect 6823 170 6857 204
rect 6823 102 6857 136
rect 6823 34 6857 68
rect 6823 -34 6857 0
rect 6823 -102 6857 -68
rect 6823 -170 6857 -136
rect 6823 -238 6857 -204
rect 6823 -306 6857 -272
rect 6823 -374 6857 -340
rect 6823 -442 6857 -408
rect 6823 -503 6857 -476
rect -277 -537 -195 -503
rect -161 -537 -127 -503
rect -93 -537 -59 -503
rect -25 -537 9 -503
rect 43 -537 77 -503
rect 111 -537 145 -503
rect 179 -537 213 -503
rect 247 -537 281 -503
rect 315 -537 349 -503
rect 383 -537 417 -503
rect 451 -537 485 -503
rect 519 -537 553 -503
rect 587 -537 621 -503
rect 655 -537 689 -503
rect 723 -537 757 -503
rect 791 -537 825 -503
rect 859 -537 893 -503
rect 927 -537 961 -503
rect 995 -537 1029 -503
rect 1063 -537 1097 -503
rect 1131 -537 1165 -503
rect 1199 -537 1233 -503
rect 1267 -537 1301 -503
rect 1335 -537 1369 -503
rect 1403 -537 1437 -503
rect 1471 -537 1505 -503
rect 1539 -537 1573 -503
rect 1607 -537 1641 -503
rect 1675 -537 1709 -503
rect 1743 -537 1777 -503
rect 1811 -537 1845 -503
rect 1879 -537 1913 -503
rect 1947 -537 1981 -503
rect 2015 -537 2049 -503
rect 2083 -537 2117 -503
rect 2151 -537 2185 -503
rect 2219 -537 2253 -503
rect 2287 -537 2321 -503
rect 2355 -537 2389 -503
rect 2423 -537 2457 -503
rect 2491 -537 2525 -503
rect 2559 -537 2593 -503
rect 2627 -537 2661 -503
rect 2695 -537 2729 -503
rect 2763 -537 2797 -503
rect 2831 -537 2865 -503
rect 2899 -537 2933 -503
rect 2967 -537 3001 -503
rect 3035 -537 3069 -503
rect 3103 -537 3137 -503
rect 3171 -537 3205 -503
rect 3239 -537 3273 -503
rect 3307 -537 3341 -503
rect 3375 -537 3409 -503
rect 3443 -537 3477 -503
rect 3511 -537 3545 -503
rect 3579 -537 3613 -503
rect 3647 -537 3681 -503
rect 3715 -537 3749 -503
rect 3783 -537 3817 -503
rect 3851 -537 3885 -503
rect 3919 -537 3953 -503
rect 3987 -537 4021 -503
rect 4055 -537 4089 -503
rect 4123 -537 4157 -503
rect 4191 -537 4225 -503
rect 4259 -537 4293 -503
rect 4327 -537 4361 -503
rect 4395 -537 4429 -503
rect 4463 -537 4497 -503
rect 4531 -537 4565 -503
rect 4599 -537 4633 -503
rect 4667 -537 4701 -503
rect 4735 -537 4769 -503
rect 4803 -537 4837 -503
rect 4871 -537 4905 -503
rect 4939 -537 4973 -503
rect 5007 -537 5041 -503
rect 5075 -537 5109 -503
rect 5143 -537 5177 -503
rect 5211 -537 5245 -503
rect 5279 -537 5313 -503
rect 5347 -537 5381 -503
rect 5415 -537 5449 -503
rect 5483 -537 5517 -503
rect 5551 -537 5585 -503
rect 5619 -537 5653 -503
rect 5687 -537 5721 -503
rect 5755 -537 5789 -503
rect 5823 -537 5857 -503
rect 5891 -537 5925 -503
rect 5959 -537 5993 -503
rect 6027 -537 6061 -503
rect 6095 -537 6129 -503
rect 6163 -537 6197 -503
rect 6231 -537 6265 -503
rect 6299 -537 6333 -503
rect 6367 -537 6401 -503
rect 6435 -537 6469 -503
rect 6503 -537 6537 -503
rect 6571 -537 6605 -503
rect 6639 -537 6673 -503
rect 6707 -537 6741 -503
rect 6775 -537 6857 -503
<< metal1 >>
rect 6467 5266 6577 5290
rect 6467 5214 6496 5266
rect 6548 5214 6577 5266
rect 60 5170 230 5210
rect 6467 5190 6577 5214
rect 57 5130 237 5170
rect 6490 5150 6570 5190
rect 60 4800 230 5130
rect 6490 5070 6660 5150
rect 60 4740 6550 4800
rect 200 4640 6550 4740
rect 60 4590 6550 4640
rect -70 4466 10 4470
rect -70 4414 -56 4466
rect -4 4414 10 4466
rect -70 4386 10 4414
rect 60 4410 250 4590
rect 370 4556 460 4560
rect 370 4504 389 4556
rect 441 4504 460 4556
rect 370 4410 460 4504
rect 670 4556 760 4560
rect 670 4504 689 4556
rect 741 4504 760 4556
rect 670 4410 760 4504
rect 970 4556 1060 4560
rect 970 4504 989 4556
rect 1041 4504 1060 4556
rect 970 4410 1060 4504
rect 1270 4556 1360 4560
rect 1270 4504 1289 4556
rect 1341 4504 1360 4556
rect 1270 4410 1360 4504
rect 1560 4466 1650 4470
rect 1560 4414 1579 4466
rect 1631 4414 1650 4466
rect 1560 4410 1650 4414
rect 1860 4466 1950 4470
rect 1860 4414 1879 4466
rect 1931 4414 1950 4466
rect 1860 4410 1950 4414
rect 2160 4466 2250 4470
rect 2160 4414 2179 4466
rect 2231 4414 2250 4466
rect 2160 4410 2250 4414
rect 2460 4466 2550 4470
rect 2460 4414 2479 4466
rect 2531 4414 2550 4466
rect 2460 4410 2550 4414
rect 2770 4466 2860 4470
rect 2770 4414 2789 4466
rect 2841 4414 2860 4466
rect 2770 4410 2860 4414
rect 3070 4466 3160 4470
rect 3070 4414 3089 4466
rect 3141 4414 3160 4466
rect 3360 4466 3550 4590
rect 5170 4556 5260 4560
rect 5170 4504 5189 4556
rect 5241 4504 5260 4556
rect 3360 4420 3389 4466
rect 3070 4410 3160 4414
rect 3370 4414 3389 4420
rect 3441 4414 3550 4466
rect 3370 4410 3550 4414
rect 3670 4466 3760 4470
rect 3670 4414 3689 4466
rect 3741 4414 3760 4466
rect 3670 4410 3760 4414
rect 3960 4466 4050 4470
rect 3960 4414 3979 4466
rect 4031 4414 4050 4466
rect 3960 4410 4050 4414
rect 4260 4466 4350 4470
rect 4260 4414 4279 4466
rect 4331 4414 4350 4466
rect 4260 4410 4350 4414
rect 4560 4466 4650 4470
rect 4560 4414 4579 4466
rect 4631 4414 4650 4466
rect 4560 4410 4650 4414
rect 4860 4466 4950 4470
rect 4860 4414 4879 4466
rect 4931 4414 4950 4466
rect 4860 4410 4950 4414
rect 5170 4410 5260 4504
rect 5470 4556 5560 4560
rect 5470 4504 5489 4556
rect 5541 4504 5560 4556
rect 5470 4410 5560 4504
rect 5770 4556 5860 4560
rect 5770 4504 5789 4556
rect 5841 4504 5860 4556
rect 5770 4410 5860 4504
rect 6070 4556 6160 4560
rect 6070 4504 6089 4556
rect 6141 4504 6160 4556
rect 6070 4410 6160 4504
rect 6360 4410 6550 4590
rect -70 4334 -56 4386
rect -4 4334 10 4386
rect -70 2226 10 4334
rect 190 2410 250 4410
rect 470 3626 550 3650
rect 470 3574 484 3626
rect 536 3574 550 3626
rect 470 3536 550 3574
rect 470 3484 484 3536
rect 536 3484 550 3536
rect 470 3446 550 3484
rect 470 3394 484 3446
rect 536 3394 550 3446
rect 470 3356 550 3394
rect 470 3304 484 3356
rect 536 3304 550 3356
rect 470 3266 550 3304
rect 470 3214 484 3266
rect 536 3214 550 3266
rect 470 3176 550 3214
rect 470 3124 484 3176
rect 536 3124 550 3176
rect 470 3110 550 3124
rect 770 3626 850 3650
rect 770 3574 784 3626
rect 836 3574 850 3626
rect 770 3536 850 3574
rect 770 3484 784 3536
rect 836 3484 850 3536
rect 770 3446 850 3484
rect 770 3394 784 3446
rect 836 3394 850 3446
rect 770 3356 850 3394
rect 770 3304 784 3356
rect 836 3304 850 3356
rect 770 3266 850 3304
rect 770 3214 784 3266
rect 836 3214 850 3266
rect 770 3176 850 3214
rect 770 3124 784 3176
rect 836 3124 850 3176
rect 770 3110 850 3124
rect 1070 3626 1150 3650
rect 1070 3574 1084 3626
rect 1136 3574 1150 3626
rect 1070 3536 1150 3574
rect 1070 3484 1084 3536
rect 1136 3484 1150 3536
rect 1070 3446 1150 3484
rect 1070 3394 1084 3446
rect 1136 3394 1150 3446
rect 1070 3356 1150 3394
rect 1070 3304 1084 3356
rect 1136 3304 1150 3356
rect 1070 3266 1150 3304
rect 1070 3214 1084 3266
rect 1136 3214 1150 3266
rect 1070 3176 1150 3214
rect 1070 3124 1084 3176
rect 1136 3124 1150 3176
rect 1070 3110 1150 3124
rect 1370 3626 1450 3650
rect 1370 3574 1384 3626
rect 1436 3574 1450 3626
rect 1370 3536 1450 3574
rect 1370 3484 1384 3536
rect 1436 3484 1450 3536
rect 1370 3446 1450 3484
rect 1370 3394 1384 3446
rect 1436 3394 1450 3446
rect 1370 3356 1450 3394
rect 1370 3304 1384 3356
rect 1436 3304 1450 3356
rect 1370 3266 1450 3304
rect 1370 3214 1384 3266
rect 1436 3214 1450 3266
rect 1370 3176 1450 3214
rect 1370 3124 1384 3176
rect 1436 3124 1450 3176
rect 1370 3110 1450 3124
rect 1670 3626 1750 3650
rect 1670 3574 1684 3626
rect 1736 3574 1750 3626
rect 1670 3536 1750 3574
rect 1670 3484 1684 3536
rect 1736 3484 1750 3536
rect 1670 3446 1750 3484
rect 1670 3394 1684 3446
rect 1736 3394 1750 3446
rect 1670 3356 1750 3394
rect 1670 3304 1684 3356
rect 1736 3304 1750 3356
rect 1670 3266 1750 3304
rect 1670 3214 1684 3266
rect 1736 3214 1750 3266
rect 1670 3176 1750 3214
rect 1670 3124 1684 3176
rect 1736 3124 1750 3176
rect 1670 3110 1750 3124
rect 1970 3626 2050 3650
rect 1970 3574 1984 3626
rect 2036 3574 2050 3626
rect 1970 3536 2050 3574
rect 1970 3484 1984 3536
rect 2036 3484 2050 3536
rect 1970 3446 2050 3484
rect 1970 3394 1984 3446
rect 2036 3394 2050 3446
rect 1970 3356 2050 3394
rect 1970 3304 1984 3356
rect 2036 3304 2050 3356
rect 1970 3266 2050 3304
rect 1970 3214 1984 3266
rect 2036 3214 2050 3266
rect 1970 3176 2050 3214
rect 1970 3124 1984 3176
rect 2036 3124 2050 3176
rect 1970 3110 2050 3124
rect 2270 3626 2350 3650
rect 2270 3574 2284 3626
rect 2336 3574 2350 3626
rect 2270 3536 2350 3574
rect 2270 3484 2284 3536
rect 2336 3484 2350 3536
rect 2270 3446 2350 3484
rect 2270 3394 2284 3446
rect 2336 3394 2350 3446
rect 2270 3356 2350 3394
rect 2270 3304 2284 3356
rect 2336 3304 2350 3356
rect 2270 3266 2350 3304
rect 2270 3214 2284 3266
rect 2336 3214 2350 3266
rect 2270 3176 2350 3214
rect 2270 3124 2284 3176
rect 2336 3124 2350 3176
rect 2270 3110 2350 3124
rect 2570 3626 2650 3650
rect 2570 3574 2584 3626
rect 2636 3574 2650 3626
rect 2570 3536 2650 3574
rect 2570 3484 2584 3536
rect 2636 3484 2650 3536
rect 2570 3446 2650 3484
rect 2570 3394 2584 3446
rect 2636 3394 2650 3446
rect 2570 3356 2650 3394
rect 2570 3304 2584 3356
rect 2636 3304 2650 3356
rect 2570 3266 2650 3304
rect 2570 3214 2584 3266
rect 2636 3214 2650 3266
rect 2570 3176 2650 3214
rect 2570 3124 2584 3176
rect 2636 3124 2650 3176
rect 2570 3110 2650 3124
rect 2870 3626 2950 3650
rect 2870 3574 2884 3626
rect 2936 3574 2950 3626
rect 2870 3536 2950 3574
rect 2870 3484 2884 3536
rect 2936 3484 2950 3536
rect 2870 3446 2950 3484
rect 2870 3394 2884 3446
rect 2936 3394 2950 3446
rect 2870 3356 2950 3394
rect 2870 3304 2884 3356
rect 2936 3304 2950 3356
rect 2870 3266 2950 3304
rect 2870 3214 2884 3266
rect 2936 3214 2950 3266
rect 2870 3176 2950 3214
rect 2870 3124 2884 3176
rect 2936 3124 2950 3176
rect 2870 3110 2950 3124
rect 3170 3626 3250 3650
rect 3170 3574 3184 3626
rect 3236 3574 3250 3626
rect 3170 3536 3250 3574
rect 3170 3484 3184 3536
rect 3236 3484 3250 3536
rect 3170 3446 3250 3484
rect 3170 3394 3184 3446
rect 3236 3394 3250 3446
rect 3170 3356 3250 3394
rect 3170 3304 3184 3356
rect 3236 3304 3250 3356
rect 3170 3266 3250 3304
rect 3170 3214 3184 3266
rect 3236 3214 3250 3266
rect 3170 3176 3250 3214
rect 3170 3124 3184 3176
rect 3236 3124 3250 3176
rect 3170 3110 3250 3124
rect 70 2370 250 2410
rect -70 2174 -56 2226
rect -4 2174 10 2226
rect -70 2146 10 2174
rect -70 2094 -56 2146
rect -4 2094 10 2146
rect -70 2090 10 2094
rect 60 2090 250 2370
rect 360 2326 460 2420
rect 360 2274 379 2326
rect 431 2274 460 2326
rect 360 2270 460 2274
rect 660 2326 760 2420
rect 660 2274 679 2326
rect 731 2274 760 2326
rect 660 2270 760 2274
rect 960 2326 1060 2420
rect 960 2274 979 2326
rect 1031 2274 1060 2326
rect 960 2270 1060 2274
rect 1260 2326 1360 2420
rect 1570 2416 1660 2420
rect 1570 2364 1589 2416
rect 1641 2364 1660 2416
rect 1570 2360 1660 2364
rect 1870 2416 1960 2420
rect 1870 2364 1889 2416
rect 1941 2364 1960 2416
rect 1870 2360 1960 2364
rect 2170 2416 2260 2420
rect 2170 2364 2189 2416
rect 2241 2364 2260 2416
rect 2170 2360 2260 2364
rect 2470 2416 2560 2420
rect 2470 2364 2489 2416
rect 2541 2364 2560 2416
rect 2890 2410 2950 3110
rect 3190 2410 3250 3110
rect 3490 2410 3550 4410
rect 3770 3626 3850 3650
rect 3770 3574 3784 3626
rect 3836 3574 3850 3626
rect 3770 3536 3850 3574
rect 3770 3484 3784 3536
rect 3836 3484 3850 3536
rect 3770 3446 3850 3484
rect 3770 3394 3784 3446
rect 3836 3394 3850 3446
rect 3770 3356 3850 3394
rect 3770 3304 3784 3356
rect 3836 3304 3850 3356
rect 3770 3266 3850 3304
rect 3770 3214 3784 3266
rect 3836 3214 3850 3266
rect 3770 3176 3850 3214
rect 3770 3124 3784 3176
rect 3836 3124 3850 3176
rect 3770 3110 3850 3124
rect 4070 3626 4150 3650
rect 4070 3574 4084 3626
rect 4136 3574 4150 3626
rect 4070 3536 4150 3574
rect 4070 3484 4084 3536
rect 4136 3484 4150 3536
rect 4070 3446 4150 3484
rect 4070 3394 4084 3446
rect 4136 3394 4150 3446
rect 4070 3356 4150 3394
rect 4070 3304 4084 3356
rect 4136 3304 4150 3356
rect 4070 3266 4150 3304
rect 4070 3214 4084 3266
rect 4136 3214 4150 3266
rect 4070 3176 4150 3214
rect 4070 3124 4084 3176
rect 4136 3124 4150 3176
rect 4070 3110 4150 3124
rect 4370 3626 4450 3650
rect 4370 3574 4384 3626
rect 4436 3574 4450 3626
rect 4370 3536 4450 3574
rect 4370 3484 4384 3536
rect 4436 3484 4450 3536
rect 4370 3446 4450 3484
rect 4370 3394 4384 3446
rect 4436 3394 4450 3446
rect 4370 3356 4450 3394
rect 4370 3304 4384 3356
rect 4436 3304 4450 3356
rect 4370 3266 4450 3304
rect 4370 3214 4384 3266
rect 4436 3214 4450 3266
rect 4370 3176 4450 3214
rect 4370 3124 4384 3176
rect 4436 3124 4450 3176
rect 4370 3110 4450 3124
rect 4670 3626 4750 3650
rect 4670 3574 4684 3626
rect 4736 3574 4750 3626
rect 4670 3536 4750 3574
rect 4670 3484 4684 3536
rect 4736 3484 4750 3536
rect 4670 3446 4750 3484
rect 4670 3394 4684 3446
rect 4736 3394 4750 3446
rect 4670 3356 4750 3394
rect 4670 3304 4684 3356
rect 4736 3304 4750 3356
rect 4670 3266 4750 3304
rect 4670 3214 4684 3266
rect 4736 3214 4750 3266
rect 4670 3176 4750 3214
rect 4670 3124 4684 3176
rect 4736 3124 4750 3176
rect 4670 3110 4750 3124
rect 4970 3626 5050 3650
rect 4970 3574 4984 3626
rect 5036 3574 5050 3626
rect 4970 3536 5050 3574
rect 4970 3484 4984 3536
rect 5036 3484 5050 3536
rect 4970 3446 5050 3484
rect 4970 3394 4984 3446
rect 5036 3394 5050 3446
rect 4970 3356 5050 3394
rect 4970 3304 4984 3356
rect 5036 3304 5050 3356
rect 4970 3266 5050 3304
rect 4970 3214 4984 3266
rect 5036 3214 5050 3266
rect 4970 3176 5050 3214
rect 4970 3124 4984 3176
rect 5036 3124 5050 3176
rect 4970 3110 5050 3124
rect 5270 3626 5350 3650
rect 5270 3574 5284 3626
rect 5336 3574 5350 3626
rect 5270 3536 5350 3574
rect 5270 3484 5284 3536
rect 5336 3484 5350 3536
rect 5270 3446 5350 3484
rect 5270 3394 5284 3446
rect 5336 3394 5350 3446
rect 5270 3356 5350 3394
rect 5270 3304 5284 3356
rect 5336 3304 5350 3356
rect 5270 3266 5350 3304
rect 5270 3214 5284 3266
rect 5336 3214 5350 3266
rect 5270 3176 5350 3214
rect 5270 3124 5284 3176
rect 5336 3124 5350 3176
rect 5270 3110 5350 3124
rect 5570 3626 5650 3650
rect 5570 3574 5584 3626
rect 5636 3574 5650 3626
rect 5570 3536 5650 3574
rect 5570 3484 5584 3536
rect 5636 3484 5650 3536
rect 5570 3446 5650 3484
rect 5570 3394 5584 3446
rect 5636 3394 5650 3446
rect 5570 3356 5650 3394
rect 5570 3304 5584 3356
rect 5636 3304 5650 3356
rect 5570 3266 5650 3304
rect 5570 3214 5584 3266
rect 5636 3214 5650 3266
rect 5570 3176 5650 3214
rect 5570 3124 5584 3176
rect 5636 3124 5650 3176
rect 5570 3110 5650 3124
rect 5870 3626 5950 3650
rect 5870 3574 5884 3626
rect 5936 3574 5950 3626
rect 5870 3536 5950 3574
rect 5870 3484 5884 3536
rect 5936 3484 5950 3536
rect 5870 3446 5950 3484
rect 5870 3394 5884 3446
rect 5936 3394 5950 3446
rect 5870 3356 5950 3394
rect 5870 3304 5884 3356
rect 5936 3304 5950 3356
rect 5870 3266 5950 3304
rect 5870 3214 5884 3266
rect 5936 3214 5950 3266
rect 5870 3176 5950 3214
rect 5870 3124 5884 3176
rect 5936 3124 5950 3176
rect 5870 3110 5950 3124
rect 6170 3626 6250 3650
rect 6170 3574 6184 3626
rect 6236 3574 6250 3626
rect 6170 3536 6250 3574
rect 6170 3484 6184 3536
rect 6236 3484 6250 3536
rect 6170 3446 6250 3484
rect 6170 3394 6184 3446
rect 6236 3394 6250 3446
rect 6170 3356 6250 3394
rect 6170 3304 6184 3356
rect 6236 3304 6250 3356
rect 6170 3266 6250 3304
rect 6170 3214 6184 3266
rect 6236 3214 6250 3266
rect 6170 3176 6250 3214
rect 6170 3124 6184 3176
rect 6236 3124 6250 3176
rect 6170 3110 6250 3124
rect 3790 2410 3850 3110
rect 2470 2360 2560 2364
rect 2770 2360 2950 2410
rect 3070 2360 3250 2410
rect 1260 2274 1279 2326
rect 1331 2274 1360 2326
rect 1260 2270 1360 2274
rect 1560 2236 1660 2240
rect 1560 2184 1589 2236
rect 1641 2184 1660 2236
rect 360 2146 450 2150
rect 360 2094 379 2146
rect 431 2094 450 2146
rect 360 2090 450 2094
rect 660 2146 750 2150
rect 660 2094 679 2146
rect 731 2094 750 2146
rect 660 2090 750 2094
rect 960 2146 1050 2150
rect 960 2094 979 2146
rect 1031 2094 1050 2146
rect 960 2090 1050 2094
rect 1260 2146 1350 2150
rect 1260 2094 1279 2146
rect 1331 2094 1350 2146
rect 1260 2090 1350 2094
rect 1560 2090 1660 2184
rect 1860 2236 1960 2240
rect 1860 2184 1889 2236
rect 1941 2184 1960 2236
rect 1860 2090 1960 2184
rect 2160 2236 2260 2240
rect 2160 2184 2189 2236
rect 2241 2184 2260 2236
rect 2160 2090 2260 2184
rect 2460 2236 2560 2240
rect 2460 2184 2489 2236
rect 2541 2184 2560 2236
rect 2460 2090 2560 2184
rect 2770 2146 2860 2150
rect 2770 2094 2789 2146
rect 2841 2094 2860 2146
rect 2770 2090 2860 2094
rect 3070 2146 3250 2150
rect 3070 2094 3089 2146
rect 3141 2094 3250 2146
rect 3070 2090 3250 2094
rect 3360 2146 3550 2410
rect 3670 2360 3850 2410
rect 3970 2416 4060 2420
rect 3970 2364 3989 2416
rect 4041 2364 4060 2416
rect 3970 2360 4060 2364
rect 4270 2416 4360 2420
rect 4270 2364 4289 2416
rect 4341 2364 4360 2416
rect 4270 2360 4360 2364
rect 4570 2416 4660 2420
rect 4570 2364 4589 2416
rect 4641 2364 4660 2416
rect 4570 2360 4660 2364
rect 4870 2416 4960 2420
rect 4870 2364 4889 2416
rect 4941 2364 4960 2416
rect 4870 2360 4960 2364
rect 5170 2326 5260 2420
rect 5170 2274 5189 2326
rect 5241 2274 5260 2326
rect 5170 2270 5260 2274
rect 5460 2326 5560 2420
rect 5460 2274 5489 2326
rect 5541 2274 5560 2326
rect 5460 2270 5560 2274
rect 5760 2326 5860 2420
rect 5760 2274 5789 2326
rect 5841 2274 5860 2326
rect 5760 2270 5860 2274
rect 6060 2326 6160 2420
rect 6490 2410 6550 4410
rect 6370 2370 6550 2410
rect 6060 2274 6089 2326
rect 6141 2274 6160 2326
rect 6060 2270 6160 2274
rect 6360 2360 6550 2370
rect 6580 4636 6660 5070
rect 6580 4584 6594 4636
rect 6646 4584 6660 4636
rect 6580 4556 6660 4584
rect 6580 4504 6594 4556
rect 6646 4504 6660 4556
rect 3960 2236 4060 2240
rect 3960 2184 3989 2236
rect 4041 2184 4060 2236
rect 3360 2094 3389 2146
rect 3441 2094 3550 2146
rect 3360 2090 3550 2094
rect 3670 2146 3760 2150
rect 3670 2094 3689 2146
rect 3741 2094 3760 2146
rect 3670 2090 3760 2094
rect 3960 2090 4060 2184
rect 4260 2236 4360 2240
rect 4260 2184 4289 2236
rect 4341 2184 4360 2236
rect 4260 2090 4360 2184
rect 4560 2236 4660 2240
rect 4560 2184 4589 2236
rect 4641 2184 4660 2236
rect 4560 2090 4660 2184
rect 4860 2236 4960 2240
rect 4860 2184 4889 2236
rect 4941 2184 4960 2236
rect 4860 2090 4960 2184
rect 6360 2150 6460 2360
rect 6580 2240 6660 4504
rect 6500 2236 6660 2240
rect 6500 2184 6514 2236
rect 6566 2184 6594 2236
rect 6646 2184 6660 2236
rect 6500 2180 6660 2184
rect 6710 4466 6790 4470
rect 6710 4414 6724 4466
rect 6776 4414 6790 4466
rect 6710 4386 6790 4414
rect 6710 4334 6724 4386
rect 6776 4334 6790 4386
rect 6710 2150 6790 4334
rect 5170 2146 5260 2150
rect 5170 2094 5189 2146
rect 5241 2094 5260 2146
rect 5170 2090 5260 2094
rect 5470 2146 5560 2150
rect 5470 2094 5489 2146
rect 5541 2094 5560 2146
rect 5470 2090 5560 2094
rect 5770 2146 5860 2150
rect 5770 2094 5789 2146
rect 5841 2094 5860 2146
rect 5770 2090 5860 2094
rect 6070 2146 6160 2150
rect 6070 2094 6089 2146
rect 6141 2094 6160 2146
rect 6070 2090 6160 2094
rect 6360 2100 6550 2150
rect 6360 2090 6460 2100
rect 190 90 250 2090
rect 470 1316 550 1340
rect 470 1264 484 1316
rect 536 1264 550 1316
rect 470 1226 550 1264
rect 470 1174 484 1226
rect 536 1174 550 1226
rect 470 1136 550 1174
rect 470 1084 484 1136
rect 536 1084 550 1136
rect 470 1046 550 1084
rect 470 994 484 1046
rect 536 994 550 1046
rect 470 956 550 994
rect 470 904 484 956
rect 536 904 550 956
rect 470 866 550 904
rect 470 814 484 866
rect 536 814 550 866
rect 470 800 550 814
rect 770 1316 850 1340
rect 770 1264 784 1316
rect 836 1264 850 1316
rect 770 1226 850 1264
rect 770 1174 784 1226
rect 836 1174 850 1226
rect 770 1136 850 1174
rect 770 1084 784 1136
rect 836 1084 850 1136
rect 770 1046 850 1084
rect 770 994 784 1046
rect 836 994 850 1046
rect 770 956 850 994
rect 770 904 784 956
rect 836 904 850 956
rect 770 866 850 904
rect 770 814 784 866
rect 836 814 850 866
rect 770 800 850 814
rect 1070 1316 1150 1340
rect 1070 1264 1084 1316
rect 1136 1264 1150 1316
rect 1070 1226 1150 1264
rect 1070 1174 1084 1226
rect 1136 1174 1150 1226
rect 1070 1136 1150 1174
rect 1070 1084 1084 1136
rect 1136 1084 1150 1136
rect 1070 1046 1150 1084
rect 1070 994 1084 1046
rect 1136 994 1150 1046
rect 1070 956 1150 994
rect 1070 904 1084 956
rect 1136 904 1150 956
rect 1070 866 1150 904
rect 1070 814 1084 866
rect 1136 814 1150 866
rect 1070 800 1150 814
rect 1370 1316 1450 1340
rect 1370 1264 1384 1316
rect 1436 1264 1450 1316
rect 1370 1226 1450 1264
rect 1370 1174 1384 1226
rect 1436 1174 1450 1226
rect 1370 1136 1450 1174
rect 1370 1084 1384 1136
rect 1436 1084 1450 1136
rect 1370 1046 1450 1084
rect 1370 994 1384 1046
rect 1436 994 1450 1046
rect 1370 956 1450 994
rect 1370 904 1384 956
rect 1436 904 1450 956
rect 1370 866 1450 904
rect 1370 814 1384 866
rect 1436 814 1450 866
rect 1370 800 1450 814
rect 1670 1316 1750 1340
rect 1670 1264 1684 1316
rect 1736 1264 1750 1316
rect 1670 1226 1750 1264
rect 1670 1174 1684 1226
rect 1736 1174 1750 1226
rect 1670 1136 1750 1174
rect 1670 1084 1684 1136
rect 1736 1084 1750 1136
rect 1670 1046 1750 1084
rect 1670 994 1684 1046
rect 1736 994 1750 1046
rect 1670 956 1750 994
rect 1670 904 1684 956
rect 1736 904 1750 956
rect 1670 866 1750 904
rect 1670 814 1684 866
rect 1736 814 1750 866
rect 1670 800 1750 814
rect 1970 1316 2050 1340
rect 1970 1264 1984 1316
rect 2036 1264 2050 1316
rect 1970 1226 2050 1264
rect 1970 1174 1984 1226
rect 2036 1174 2050 1226
rect 1970 1136 2050 1174
rect 1970 1084 1984 1136
rect 2036 1084 2050 1136
rect 1970 1046 2050 1084
rect 1970 994 1984 1046
rect 2036 994 2050 1046
rect 1970 956 2050 994
rect 1970 904 1984 956
rect 2036 904 2050 956
rect 1970 866 2050 904
rect 1970 814 1984 866
rect 2036 814 2050 866
rect 1970 800 2050 814
rect 2270 1316 2350 1340
rect 2270 1264 2284 1316
rect 2336 1264 2350 1316
rect 2270 1226 2350 1264
rect 2270 1174 2284 1226
rect 2336 1174 2350 1226
rect 2270 1136 2350 1174
rect 2270 1084 2284 1136
rect 2336 1084 2350 1136
rect 2270 1046 2350 1084
rect 2270 994 2284 1046
rect 2336 994 2350 1046
rect 2270 956 2350 994
rect 2270 904 2284 956
rect 2336 904 2350 956
rect 2270 866 2350 904
rect 2270 814 2284 866
rect 2336 814 2350 866
rect 2270 800 2350 814
rect 2570 1316 2650 1340
rect 2570 1264 2584 1316
rect 2636 1264 2650 1316
rect 2570 1226 2650 1264
rect 2570 1174 2584 1226
rect 2636 1174 2650 1226
rect 2570 1136 2650 1174
rect 2570 1084 2584 1136
rect 2636 1084 2650 1136
rect 2570 1046 2650 1084
rect 2570 994 2584 1046
rect 2636 994 2650 1046
rect 2570 956 2650 994
rect 2570 904 2584 956
rect 2636 904 2650 956
rect 2570 866 2650 904
rect 2570 814 2584 866
rect 2636 814 2650 866
rect 2570 800 2650 814
rect 2870 1316 2950 1340
rect 2870 1264 2884 1316
rect 2936 1264 2950 1316
rect 2870 1226 2950 1264
rect 2870 1174 2884 1226
rect 2936 1174 2950 1226
rect 2870 1136 2950 1174
rect 2870 1084 2884 1136
rect 2936 1084 2950 1136
rect 2870 1046 2950 1084
rect 2870 994 2884 1046
rect 2936 994 2950 1046
rect 2870 956 2950 994
rect 2870 904 2884 956
rect 2936 904 2950 956
rect 2870 866 2950 904
rect 2870 814 2884 866
rect 2936 814 2950 866
rect 2870 800 2950 814
rect 2890 100 2950 800
rect 60 -80 250 90
rect 360 96 450 100
rect 360 44 379 96
rect 431 44 450 96
rect 360 40 450 44
rect 660 96 750 100
rect 660 44 679 96
rect 731 44 750 96
rect 660 40 750 44
rect 960 96 1050 100
rect 960 44 979 96
rect 1031 44 1050 96
rect 960 40 1050 44
rect 1260 96 1350 100
rect 1260 44 1279 96
rect 1331 44 1350 96
rect 1260 40 1350 44
rect 1560 6 1660 90
rect 1560 -46 1579 6
rect 1631 -46 1660 6
rect 1560 -50 1660 -46
rect 1860 6 1960 90
rect 1860 -46 1879 6
rect 1931 -46 1960 6
rect 1860 -50 1960 -46
rect 2160 6 2260 90
rect 2160 -46 2179 6
rect 2231 -46 2260 6
rect 2160 -50 2260 -46
rect 2460 6 2560 90
rect 2770 40 2950 100
rect 3190 90 3250 2090
rect 3470 1316 3550 1340
rect 3470 1264 3484 1316
rect 3536 1264 3550 1316
rect 3470 1226 3550 1264
rect 3470 1174 3484 1226
rect 3536 1174 3550 1226
rect 3470 1136 3550 1174
rect 3470 1084 3484 1136
rect 3536 1084 3550 1136
rect 3470 1046 3550 1084
rect 3470 994 3484 1046
rect 3536 994 3550 1046
rect 3470 956 3550 994
rect 3470 904 3484 956
rect 3536 904 3550 956
rect 3470 866 3550 904
rect 3470 814 3484 866
rect 3536 814 3550 866
rect 3470 800 3550 814
rect 3770 1316 3850 1340
rect 3770 1264 3784 1316
rect 3836 1264 3850 1316
rect 3770 1226 3850 1264
rect 3770 1174 3784 1226
rect 3836 1174 3850 1226
rect 3770 1136 3850 1174
rect 3770 1084 3784 1136
rect 3836 1084 3850 1136
rect 3770 1046 3850 1084
rect 3770 994 3784 1046
rect 3836 994 3850 1046
rect 3770 956 3850 994
rect 3770 904 3784 956
rect 3836 904 3850 956
rect 3770 866 3850 904
rect 3770 814 3784 866
rect 3836 814 3850 866
rect 3770 800 3850 814
rect 4070 1316 4150 1340
rect 4070 1264 4084 1316
rect 4136 1264 4150 1316
rect 4070 1226 4150 1264
rect 4070 1174 4084 1226
rect 4136 1174 4150 1226
rect 4070 1136 4150 1174
rect 4070 1084 4084 1136
rect 4136 1084 4150 1136
rect 4070 1046 4150 1084
rect 4070 994 4084 1046
rect 4136 994 4150 1046
rect 4070 956 4150 994
rect 4070 904 4084 956
rect 4136 904 4150 956
rect 4070 866 4150 904
rect 4070 814 4084 866
rect 4136 814 4150 866
rect 4070 800 4150 814
rect 4370 1316 4450 1340
rect 4370 1264 4384 1316
rect 4436 1264 4450 1316
rect 4370 1226 4450 1264
rect 4370 1174 4384 1226
rect 4436 1174 4450 1226
rect 4370 1136 4450 1174
rect 4370 1084 4384 1136
rect 4436 1084 4450 1136
rect 4370 1046 4450 1084
rect 4370 994 4384 1046
rect 4436 994 4450 1046
rect 4370 956 4450 994
rect 4370 904 4384 956
rect 4436 904 4450 956
rect 4370 866 4450 904
rect 4370 814 4384 866
rect 4436 814 4450 866
rect 4370 800 4450 814
rect 4670 1316 4750 1340
rect 4670 1264 4684 1316
rect 4736 1264 4750 1316
rect 4670 1226 4750 1264
rect 4670 1174 4684 1226
rect 4736 1174 4750 1226
rect 4670 1136 4750 1174
rect 4670 1084 4684 1136
rect 4736 1084 4750 1136
rect 4670 1046 4750 1084
rect 4670 994 4684 1046
rect 4736 994 4750 1046
rect 4670 956 4750 994
rect 4670 904 4684 956
rect 4736 904 4750 956
rect 4670 866 4750 904
rect 4670 814 4684 866
rect 4736 814 4750 866
rect 4670 800 4750 814
rect 4970 1316 5050 1340
rect 4970 1264 4984 1316
rect 5036 1264 5050 1316
rect 4970 1226 5050 1264
rect 4970 1174 4984 1226
rect 5036 1174 5050 1226
rect 4970 1136 5050 1174
rect 4970 1084 4984 1136
rect 5036 1084 5050 1136
rect 4970 1046 5050 1084
rect 4970 994 4984 1046
rect 5036 994 5050 1046
rect 4970 956 5050 994
rect 4970 904 4984 956
rect 5036 904 5050 956
rect 4970 866 5050 904
rect 4970 814 4984 866
rect 5036 814 5050 866
rect 4970 800 5050 814
rect 5270 1316 5350 1340
rect 5270 1264 5284 1316
rect 5336 1264 5350 1316
rect 5270 1226 5350 1264
rect 5270 1174 5284 1226
rect 5336 1174 5350 1226
rect 5270 1136 5350 1174
rect 5270 1084 5284 1136
rect 5336 1084 5350 1136
rect 5270 1046 5350 1084
rect 5270 994 5284 1046
rect 5336 994 5350 1046
rect 5270 956 5350 994
rect 5270 904 5284 956
rect 5336 904 5350 956
rect 5270 866 5350 904
rect 5270 814 5284 866
rect 5336 814 5350 866
rect 5270 800 5350 814
rect 5570 1316 5650 1340
rect 5570 1264 5584 1316
rect 5636 1264 5650 1316
rect 5570 1226 5650 1264
rect 5570 1174 5584 1226
rect 5636 1174 5650 1226
rect 5570 1136 5650 1174
rect 5570 1084 5584 1136
rect 5636 1084 5650 1136
rect 5570 1046 5650 1084
rect 5570 994 5584 1046
rect 5636 994 5650 1046
rect 5570 956 5650 994
rect 5570 904 5584 956
rect 5636 904 5650 956
rect 5570 866 5650 904
rect 5570 814 5584 866
rect 5636 814 5650 866
rect 5570 800 5650 814
rect 5870 1316 5950 1340
rect 5870 1264 5884 1316
rect 5936 1264 5950 1316
rect 5870 1226 5950 1264
rect 5870 1174 5884 1226
rect 5936 1174 5950 1226
rect 5870 1136 5950 1174
rect 5870 1084 5884 1136
rect 5936 1084 5950 1136
rect 5870 1046 5950 1084
rect 5870 994 5884 1046
rect 5936 994 5950 1046
rect 5870 956 5950 994
rect 5870 904 5884 956
rect 5936 904 5950 956
rect 5870 866 5950 904
rect 5870 814 5884 866
rect 5936 814 5950 866
rect 5870 800 5950 814
rect 6170 1316 6250 1340
rect 6170 1264 6184 1316
rect 6236 1264 6250 1316
rect 6170 1226 6250 1264
rect 6170 1174 6184 1226
rect 6236 1174 6250 1226
rect 6170 1136 6250 1174
rect 6170 1084 6184 1136
rect 6236 1084 6250 1136
rect 6170 1046 6250 1084
rect 6170 994 6184 1046
rect 6236 994 6250 1046
rect 6170 956 6250 994
rect 6170 904 6184 956
rect 6236 904 6250 956
rect 6170 866 6250 904
rect 6170 814 6184 866
rect 6236 814 6250 866
rect 6170 800 6250 814
rect 3490 100 3550 800
rect 3790 100 3850 800
rect 2460 -46 2479 6
rect 2531 -46 2560 6
rect 2460 -50 2560 -46
rect 3060 -80 3250 90
rect 3370 40 3550 100
rect 3670 40 3850 100
rect 5170 96 5260 100
rect 3970 6 4070 90
rect 3970 -46 3989 6
rect 4041 -46 4070 6
rect 3970 -50 4070 -46
rect 4260 6 4360 90
rect 4260 -46 4289 6
rect 4341 -46 4360 6
rect 4260 -50 4360 -46
rect 4560 6 4660 90
rect 4560 -46 4589 6
rect 4641 -46 4660 6
rect 4560 -50 4660 -46
rect 4860 6 4960 90
rect 5170 44 5189 96
rect 5241 44 5260 96
rect 5170 40 5260 44
rect 5470 96 5560 100
rect 5470 44 5489 96
rect 5541 44 5560 96
rect 5470 40 5560 44
rect 5770 96 5860 100
rect 5770 44 5789 96
rect 5841 44 5860 96
rect 5770 40 5860 44
rect 6070 96 6160 100
rect 6070 44 6089 96
rect 6141 44 6160 96
rect 6490 90 6550 2100
rect 6630 2146 6790 2150
rect 6630 2094 6644 2146
rect 6696 2094 6724 2146
rect 6776 2094 6790 2146
rect 6630 2090 6790 2094
rect 6070 40 6160 44
rect 4860 -46 4889 6
rect 4941 -46 4960 6
rect 4860 -50 4960 -46
rect 6360 -80 6550 90
rect 60 -130 6550 -80
rect 190 -230 6550 -130
rect 60 -290 6550 -230
<< via1 >>
rect 6496 5214 6548 5266
rect -56 4414 -4 4466
rect 389 4504 441 4556
rect 689 4504 741 4556
rect 989 4504 1041 4556
rect 1289 4504 1341 4556
rect 1579 4414 1631 4466
rect 1879 4414 1931 4466
rect 2179 4414 2231 4466
rect 2479 4414 2531 4466
rect 2789 4414 2841 4466
rect 3089 4414 3141 4466
rect 5189 4504 5241 4556
rect 3389 4414 3441 4466
rect 3689 4414 3741 4466
rect 3979 4414 4031 4466
rect 4279 4414 4331 4466
rect 4579 4414 4631 4466
rect 4879 4414 4931 4466
rect 5489 4504 5541 4556
rect 5789 4504 5841 4556
rect 6089 4504 6141 4556
rect -56 4334 -4 4386
rect 484 3574 536 3626
rect 484 3484 536 3536
rect 484 3394 536 3446
rect 484 3304 536 3356
rect 484 3214 536 3266
rect 484 3124 536 3176
rect 784 3574 836 3626
rect 784 3484 836 3536
rect 784 3394 836 3446
rect 784 3304 836 3356
rect 784 3214 836 3266
rect 784 3124 836 3176
rect 1084 3574 1136 3626
rect 1084 3484 1136 3536
rect 1084 3394 1136 3446
rect 1084 3304 1136 3356
rect 1084 3214 1136 3266
rect 1084 3124 1136 3176
rect 1384 3574 1436 3626
rect 1384 3484 1436 3536
rect 1384 3394 1436 3446
rect 1384 3304 1436 3356
rect 1384 3214 1436 3266
rect 1384 3124 1436 3176
rect 1684 3574 1736 3626
rect 1684 3484 1736 3536
rect 1684 3394 1736 3446
rect 1684 3304 1736 3356
rect 1684 3214 1736 3266
rect 1684 3124 1736 3176
rect 1984 3574 2036 3626
rect 1984 3484 2036 3536
rect 1984 3394 2036 3446
rect 1984 3304 2036 3356
rect 1984 3214 2036 3266
rect 1984 3124 2036 3176
rect 2284 3574 2336 3626
rect 2284 3484 2336 3536
rect 2284 3394 2336 3446
rect 2284 3304 2336 3356
rect 2284 3214 2336 3266
rect 2284 3124 2336 3176
rect 2584 3574 2636 3626
rect 2584 3484 2636 3536
rect 2584 3394 2636 3446
rect 2584 3304 2636 3356
rect 2584 3214 2636 3266
rect 2584 3124 2636 3176
rect 2884 3574 2936 3626
rect 2884 3484 2936 3536
rect 2884 3394 2936 3446
rect 2884 3304 2936 3356
rect 2884 3214 2936 3266
rect 2884 3124 2936 3176
rect 3184 3574 3236 3626
rect 3184 3484 3236 3536
rect 3184 3394 3236 3446
rect 3184 3304 3236 3356
rect 3184 3214 3236 3266
rect 3184 3124 3236 3176
rect -56 2174 -4 2226
rect -56 2094 -4 2146
rect 379 2274 431 2326
rect 679 2274 731 2326
rect 979 2274 1031 2326
rect 1589 2364 1641 2416
rect 1889 2364 1941 2416
rect 2189 2364 2241 2416
rect 2489 2364 2541 2416
rect 3784 3574 3836 3626
rect 3784 3484 3836 3536
rect 3784 3394 3836 3446
rect 3784 3304 3836 3356
rect 3784 3214 3836 3266
rect 3784 3124 3836 3176
rect 4084 3574 4136 3626
rect 4084 3484 4136 3536
rect 4084 3394 4136 3446
rect 4084 3304 4136 3356
rect 4084 3214 4136 3266
rect 4084 3124 4136 3176
rect 4384 3574 4436 3626
rect 4384 3484 4436 3536
rect 4384 3394 4436 3446
rect 4384 3304 4436 3356
rect 4384 3214 4436 3266
rect 4384 3124 4436 3176
rect 4684 3574 4736 3626
rect 4684 3484 4736 3536
rect 4684 3394 4736 3446
rect 4684 3304 4736 3356
rect 4684 3214 4736 3266
rect 4684 3124 4736 3176
rect 4984 3574 5036 3626
rect 4984 3484 5036 3536
rect 4984 3394 5036 3446
rect 4984 3304 5036 3356
rect 4984 3214 5036 3266
rect 4984 3124 5036 3176
rect 5284 3574 5336 3626
rect 5284 3484 5336 3536
rect 5284 3394 5336 3446
rect 5284 3304 5336 3356
rect 5284 3214 5336 3266
rect 5284 3124 5336 3176
rect 5584 3574 5636 3626
rect 5584 3484 5636 3536
rect 5584 3394 5636 3446
rect 5584 3304 5636 3356
rect 5584 3214 5636 3266
rect 5584 3124 5636 3176
rect 5884 3574 5936 3626
rect 5884 3484 5936 3536
rect 5884 3394 5936 3446
rect 5884 3304 5936 3356
rect 5884 3214 5936 3266
rect 5884 3124 5936 3176
rect 6184 3574 6236 3626
rect 6184 3484 6236 3536
rect 6184 3394 6236 3446
rect 6184 3304 6236 3356
rect 6184 3214 6236 3266
rect 6184 3124 6236 3176
rect 1279 2274 1331 2326
rect 1589 2184 1641 2236
rect 379 2094 431 2146
rect 679 2094 731 2146
rect 979 2094 1031 2146
rect 1279 2094 1331 2146
rect 1889 2184 1941 2236
rect 2189 2184 2241 2236
rect 2489 2184 2541 2236
rect 2789 2094 2841 2146
rect 3089 2094 3141 2146
rect 3989 2364 4041 2416
rect 4289 2364 4341 2416
rect 4589 2364 4641 2416
rect 4889 2364 4941 2416
rect 5189 2274 5241 2326
rect 5489 2274 5541 2326
rect 5789 2274 5841 2326
rect 6089 2274 6141 2326
rect 6594 4584 6646 4636
rect 6594 4504 6646 4556
rect 3989 2184 4041 2236
rect 3389 2094 3441 2146
rect 3689 2094 3741 2146
rect 4289 2184 4341 2236
rect 4589 2184 4641 2236
rect 4889 2184 4941 2236
rect 6514 2184 6566 2236
rect 6594 2184 6646 2236
rect 6724 4414 6776 4466
rect 6724 4334 6776 4386
rect 5189 2094 5241 2146
rect 5489 2094 5541 2146
rect 5789 2094 5841 2146
rect 6089 2094 6141 2146
rect 484 1264 536 1316
rect 484 1174 536 1226
rect 484 1084 536 1136
rect 484 994 536 1046
rect 484 904 536 956
rect 484 814 536 866
rect 784 1264 836 1316
rect 784 1174 836 1226
rect 784 1084 836 1136
rect 784 994 836 1046
rect 784 904 836 956
rect 784 814 836 866
rect 1084 1264 1136 1316
rect 1084 1174 1136 1226
rect 1084 1084 1136 1136
rect 1084 994 1136 1046
rect 1084 904 1136 956
rect 1084 814 1136 866
rect 1384 1264 1436 1316
rect 1384 1174 1436 1226
rect 1384 1084 1436 1136
rect 1384 994 1436 1046
rect 1384 904 1436 956
rect 1384 814 1436 866
rect 1684 1264 1736 1316
rect 1684 1174 1736 1226
rect 1684 1084 1736 1136
rect 1684 994 1736 1046
rect 1684 904 1736 956
rect 1684 814 1736 866
rect 1984 1264 2036 1316
rect 1984 1174 2036 1226
rect 1984 1084 2036 1136
rect 1984 994 2036 1046
rect 1984 904 2036 956
rect 1984 814 2036 866
rect 2284 1264 2336 1316
rect 2284 1174 2336 1226
rect 2284 1084 2336 1136
rect 2284 994 2336 1046
rect 2284 904 2336 956
rect 2284 814 2336 866
rect 2584 1264 2636 1316
rect 2584 1174 2636 1226
rect 2584 1084 2636 1136
rect 2584 994 2636 1046
rect 2584 904 2636 956
rect 2584 814 2636 866
rect 2884 1264 2936 1316
rect 2884 1174 2936 1226
rect 2884 1084 2936 1136
rect 2884 994 2936 1046
rect 2884 904 2936 956
rect 2884 814 2936 866
rect 379 44 431 96
rect 679 44 731 96
rect 979 44 1031 96
rect 1279 44 1331 96
rect 1579 -46 1631 6
rect 1879 -46 1931 6
rect 2179 -46 2231 6
rect 3484 1264 3536 1316
rect 3484 1174 3536 1226
rect 3484 1084 3536 1136
rect 3484 994 3536 1046
rect 3484 904 3536 956
rect 3484 814 3536 866
rect 3784 1264 3836 1316
rect 3784 1174 3836 1226
rect 3784 1084 3836 1136
rect 3784 994 3836 1046
rect 3784 904 3836 956
rect 3784 814 3836 866
rect 4084 1264 4136 1316
rect 4084 1174 4136 1226
rect 4084 1084 4136 1136
rect 4084 994 4136 1046
rect 4084 904 4136 956
rect 4084 814 4136 866
rect 4384 1264 4436 1316
rect 4384 1174 4436 1226
rect 4384 1084 4436 1136
rect 4384 994 4436 1046
rect 4384 904 4436 956
rect 4384 814 4436 866
rect 4684 1264 4736 1316
rect 4684 1174 4736 1226
rect 4684 1084 4736 1136
rect 4684 994 4736 1046
rect 4684 904 4736 956
rect 4684 814 4736 866
rect 4984 1264 5036 1316
rect 4984 1174 5036 1226
rect 4984 1084 5036 1136
rect 4984 994 5036 1046
rect 4984 904 5036 956
rect 4984 814 5036 866
rect 5284 1264 5336 1316
rect 5284 1174 5336 1226
rect 5284 1084 5336 1136
rect 5284 994 5336 1046
rect 5284 904 5336 956
rect 5284 814 5336 866
rect 5584 1264 5636 1316
rect 5584 1174 5636 1226
rect 5584 1084 5636 1136
rect 5584 994 5636 1046
rect 5584 904 5636 956
rect 5584 814 5636 866
rect 5884 1264 5936 1316
rect 5884 1174 5936 1226
rect 5884 1084 5936 1136
rect 5884 994 5936 1046
rect 5884 904 5936 956
rect 5884 814 5936 866
rect 6184 1264 6236 1316
rect 6184 1174 6236 1226
rect 6184 1084 6236 1136
rect 6184 994 6236 1046
rect 6184 904 6236 956
rect 6184 814 6236 866
rect 2479 -46 2531 6
rect 3989 -46 4041 6
rect 4289 -46 4341 6
rect 4589 -46 4641 6
rect 5189 44 5241 96
rect 5489 44 5541 96
rect 5789 44 5841 96
rect 6089 44 6141 96
rect 6644 2094 6696 2146
rect 6724 2094 6776 2146
rect 4889 -46 4941 6
<< metal2 >>
rect 6467 5268 6577 5290
rect 6467 5212 6494 5268
rect 6550 5212 6577 5268
rect 6467 5190 6577 5212
rect 6707 5268 6817 5290
rect 6707 5212 6734 5268
rect 6790 5212 6817 5268
rect 6707 5190 6817 5212
rect 6710 4890 6790 5190
rect -70 4830 6790 4890
rect -70 4470 10 4830
rect 6580 4636 6660 4640
rect 6580 4584 6594 4636
rect 6646 4584 6660 4636
rect 6580 4560 6660 4584
rect 370 4556 6660 4560
rect 370 4504 389 4556
rect 441 4504 689 4556
rect 741 4504 989 4556
rect 1041 4504 1289 4556
rect 1341 4504 5189 4556
rect 5241 4504 5489 4556
rect 5541 4504 5789 4556
rect 5841 4504 6089 4556
rect 6141 4504 6594 4556
rect 6646 4504 6660 4556
rect 370 4500 6660 4504
rect 6710 4470 6790 4830
rect -70 4466 2550 4470
rect -70 4414 -56 4466
rect -4 4414 1579 4466
rect 1631 4414 1879 4466
rect 1931 4414 2179 4466
rect 2231 4414 2479 4466
rect 2531 4414 2550 4466
rect -70 4410 2550 4414
rect 2770 4466 3760 4470
rect 2770 4414 2789 4466
rect 2841 4414 3089 4466
rect 3141 4414 3389 4466
rect 3441 4414 3689 4466
rect 3741 4414 3760 4466
rect 2770 4410 3760 4414
rect 3960 4466 6790 4470
rect 3960 4414 3979 4466
rect 4031 4414 4279 4466
rect 4331 4414 4579 4466
rect 4631 4414 4879 4466
rect 4931 4414 6724 4466
rect 6776 4414 6790 4466
rect 3960 4410 6790 4414
rect -70 4386 10 4410
rect -70 4334 -56 4386
rect -4 4334 10 4386
rect -70 4330 10 4334
rect 6710 4386 6790 4410
rect 6710 4334 6724 4386
rect 6776 4334 6790 4386
rect 6710 4330 6790 4334
rect 470 3628 550 3650
rect 470 3572 482 3628
rect 538 3572 550 3628
rect 470 3538 550 3572
rect 470 3482 482 3538
rect 538 3482 550 3538
rect 470 3448 550 3482
rect 470 3392 482 3448
rect 538 3392 550 3448
rect 470 3358 550 3392
rect 470 3302 482 3358
rect 538 3302 550 3358
rect 470 3268 550 3302
rect 470 3212 482 3268
rect 538 3212 550 3268
rect 470 3178 550 3212
rect 470 3122 482 3178
rect 538 3122 550 3178
rect 470 3110 550 3122
rect 770 3628 850 3650
rect 770 3572 782 3628
rect 838 3572 850 3628
rect 770 3538 850 3572
rect 770 3482 782 3538
rect 838 3482 850 3538
rect 770 3448 850 3482
rect 770 3392 782 3448
rect 838 3392 850 3448
rect 770 3358 850 3392
rect 770 3302 782 3358
rect 838 3302 850 3358
rect 770 3268 850 3302
rect 770 3212 782 3268
rect 838 3212 850 3268
rect 770 3178 850 3212
rect 770 3122 782 3178
rect 838 3122 850 3178
rect 770 3110 850 3122
rect 1070 3628 1150 3650
rect 1070 3572 1082 3628
rect 1138 3572 1150 3628
rect 1070 3538 1150 3572
rect 1070 3482 1082 3538
rect 1138 3482 1150 3538
rect 1070 3448 1150 3482
rect 1070 3392 1082 3448
rect 1138 3392 1150 3448
rect 1070 3358 1150 3392
rect 1070 3302 1082 3358
rect 1138 3302 1150 3358
rect 1070 3268 1150 3302
rect 1070 3212 1082 3268
rect 1138 3212 1150 3268
rect 1070 3178 1150 3212
rect 1070 3122 1082 3178
rect 1138 3122 1150 3178
rect 1070 3110 1150 3122
rect 1370 3628 1450 3650
rect 1370 3572 1382 3628
rect 1438 3572 1450 3628
rect 1370 3538 1450 3572
rect 1370 3482 1382 3538
rect 1438 3482 1450 3538
rect 1370 3448 1450 3482
rect 1370 3392 1382 3448
rect 1438 3392 1450 3448
rect 1370 3358 1450 3392
rect 1370 3302 1382 3358
rect 1438 3302 1450 3358
rect 1370 3268 1450 3302
rect 1370 3212 1382 3268
rect 1438 3212 1450 3268
rect 1370 3178 1450 3212
rect 1370 3122 1382 3178
rect 1438 3122 1450 3178
rect 1370 3110 1450 3122
rect 1670 3628 1750 3650
rect 1670 3572 1682 3628
rect 1738 3572 1750 3628
rect 1670 3538 1750 3572
rect 1670 3482 1682 3538
rect 1738 3482 1750 3538
rect 1670 3448 1750 3482
rect 1670 3392 1682 3448
rect 1738 3392 1750 3448
rect 1670 3358 1750 3392
rect 1670 3302 1682 3358
rect 1738 3302 1750 3358
rect 1670 3268 1750 3302
rect 1670 3212 1682 3268
rect 1738 3212 1750 3268
rect 1670 3178 1750 3212
rect 1670 3122 1682 3178
rect 1738 3122 1750 3178
rect 1670 3110 1750 3122
rect 1970 3628 2050 3650
rect 1970 3572 1982 3628
rect 2038 3572 2050 3628
rect 1970 3538 2050 3572
rect 1970 3482 1982 3538
rect 2038 3482 2050 3538
rect 1970 3448 2050 3482
rect 1970 3392 1982 3448
rect 2038 3392 2050 3448
rect 1970 3358 2050 3392
rect 1970 3302 1982 3358
rect 2038 3302 2050 3358
rect 1970 3268 2050 3302
rect 1970 3212 1982 3268
rect 2038 3212 2050 3268
rect 1970 3178 2050 3212
rect 1970 3122 1982 3178
rect 2038 3122 2050 3178
rect 1970 3110 2050 3122
rect 2270 3628 2350 3650
rect 2270 3572 2282 3628
rect 2338 3572 2350 3628
rect 2270 3538 2350 3572
rect 2270 3482 2282 3538
rect 2338 3482 2350 3538
rect 2270 3448 2350 3482
rect 2270 3392 2282 3448
rect 2338 3392 2350 3448
rect 2270 3358 2350 3392
rect 2270 3302 2282 3358
rect 2338 3302 2350 3358
rect 2270 3268 2350 3302
rect 2270 3212 2282 3268
rect 2338 3212 2350 3268
rect 2270 3178 2350 3212
rect 2270 3122 2282 3178
rect 2338 3122 2350 3178
rect 2270 3110 2350 3122
rect 2570 3628 2650 3650
rect 2570 3572 2582 3628
rect 2638 3572 2650 3628
rect 2570 3538 2650 3572
rect 2570 3482 2582 3538
rect 2638 3482 2650 3538
rect 2570 3448 2650 3482
rect 2570 3392 2582 3448
rect 2638 3392 2650 3448
rect 2570 3358 2650 3392
rect 2570 3302 2582 3358
rect 2638 3302 2650 3358
rect 2570 3268 2650 3302
rect 2570 3212 2582 3268
rect 2638 3212 2650 3268
rect 2570 3178 2650 3212
rect 2570 3122 2582 3178
rect 2638 3122 2650 3178
rect 2570 3110 2650 3122
rect 2870 3628 2950 3650
rect 2870 3572 2882 3628
rect 2938 3572 2950 3628
rect 2870 3538 2950 3572
rect 2870 3482 2882 3538
rect 2938 3482 2950 3538
rect 2870 3448 2950 3482
rect 2870 3392 2882 3448
rect 2938 3392 2950 3448
rect 2870 3358 2950 3392
rect 2870 3302 2882 3358
rect 2938 3302 2950 3358
rect 2870 3268 2950 3302
rect 2870 3212 2882 3268
rect 2938 3212 2950 3268
rect 2870 3178 2950 3212
rect 2870 3122 2882 3178
rect 2938 3122 2950 3178
rect 2870 3110 2950 3122
rect 3170 3628 3250 3650
rect 3170 3572 3182 3628
rect 3238 3572 3250 3628
rect 3170 3538 3250 3572
rect 3170 3482 3182 3538
rect 3238 3482 3250 3538
rect 3170 3448 3250 3482
rect 3170 3392 3182 3448
rect 3238 3392 3250 3448
rect 3170 3358 3250 3392
rect 3170 3302 3182 3358
rect 3238 3302 3250 3358
rect 3170 3268 3250 3302
rect 3170 3212 3182 3268
rect 3238 3212 3250 3268
rect 3170 3178 3250 3212
rect 3170 3122 3182 3178
rect 3238 3122 3250 3178
rect 3170 3110 3250 3122
rect 3770 3628 3850 3650
rect 3770 3572 3782 3628
rect 3838 3572 3850 3628
rect 3770 3538 3850 3572
rect 3770 3482 3782 3538
rect 3838 3482 3850 3538
rect 3770 3448 3850 3482
rect 3770 3392 3782 3448
rect 3838 3392 3850 3448
rect 3770 3358 3850 3392
rect 3770 3302 3782 3358
rect 3838 3302 3850 3358
rect 3770 3268 3850 3302
rect 3770 3212 3782 3268
rect 3838 3212 3850 3268
rect 3770 3178 3850 3212
rect 3770 3122 3782 3178
rect 3838 3122 3850 3178
rect 3770 3110 3850 3122
rect 4070 3628 4150 3650
rect 4070 3572 4082 3628
rect 4138 3572 4150 3628
rect 4070 3538 4150 3572
rect 4070 3482 4082 3538
rect 4138 3482 4150 3538
rect 4070 3448 4150 3482
rect 4070 3392 4082 3448
rect 4138 3392 4150 3448
rect 4070 3358 4150 3392
rect 4070 3302 4082 3358
rect 4138 3302 4150 3358
rect 4070 3268 4150 3302
rect 4070 3212 4082 3268
rect 4138 3212 4150 3268
rect 4070 3178 4150 3212
rect 4070 3122 4082 3178
rect 4138 3122 4150 3178
rect 4070 3110 4150 3122
rect 4370 3628 4450 3650
rect 4370 3572 4382 3628
rect 4438 3572 4450 3628
rect 4370 3538 4450 3572
rect 4370 3482 4382 3538
rect 4438 3482 4450 3538
rect 4370 3448 4450 3482
rect 4370 3392 4382 3448
rect 4438 3392 4450 3448
rect 4370 3358 4450 3392
rect 4370 3302 4382 3358
rect 4438 3302 4450 3358
rect 4370 3268 4450 3302
rect 4370 3212 4382 3268
rect 4438 3212 4450 3268
rect 4370 3178 4450 3212
rect 4370 3122 4382 3178
rect 4438 3122 4450 3178
rect 4370 3110 4450 3122
rect 4670 3628 4750 3650
rect 4670 3572 4682 3628
rect 4738 3572 4750 3628
rect 4670 3538 4750 3572
rect 4670 3482 4682 3538
rect 4738 3482 4750 3538
rect 4670 3448 4750 3482
rect 4670 3392 4682 3448
rect 4738 3392 4750 3448
rect 4670 3358 4750 3392
rect 4670 3302 4682 3358
rect 4738 3302 4750 3358
rect 4670 3268 4750 3302
rect 4670 3212 4682 3268
rect 4738 3212 4750 3268
rect 4670 3178 4750 3212
rect 4670 3122 4682 3178
rect 4738 3122 4750 3178
rect 4670 3110 4750 3122
rect 4970 3628 5050 3650
rect 4970 3572 4982 3628
rect 5038 3572 5050 3628
rect 4970 3538 5050 3572
rect 4970 3482 4982 3538
rect 5038 3482 5050 3538
rect 4970 3448 5050 3482
rect 4970 3392 4982 3448
rect 5038 3392 5050 3448
rect 4970 3358 5050 3392
rect 4970 3302 4982 3358
rect 5038 3302 5050 3358
rect 4970 3268 5050 3302
rect 4970 3212 4982 3268
rect 5038 3212 5050 3268
rect 4970 3178 5050 3212
rect 4970 3122 4982 3178
rect 5038 3122 5050 3178
rect 4970 3110 5050 3122
rect 5270 3628 5350 3650
rect 5270 3572 5282 3628
rect 5338 3572 5350 3628
rect 5270 3538 5350 3572
rect 5270 3482 5282 3538
rect 5338 3482 5350 3538
rect 5270 3448 5350 3482
rect 5270 3392 5282 3448
rect 5338 3392 5350 3448
rect 5270 3358 5350 3392
rect 5270 3302 5282 3358
rect 5338 3302 5350 3358
rect 5270 3268 5350 3302
rect 5270 3212 5282 3268
rect 5338 3212 5350 3268
rect 5270 3178 5350 3212
rect 5270 3122 5282 3178
rect 5338 3122 5350 3178
rect 5270 3110 5350 3122
rect 5570 3628 5650 3650
rect 5570 3572 5582 3628
rect 5638 3572 5650 3628
rect 5570 3538 5650 3572
rect 5570 3482 5582 3538
rect 5638 3482 5650 3538
rect 5570 3448 5650 3482
rect 5570 3392 5582 3448
rect 5638 3392 5650 3448
rect 5570 3358 5650 3392
rect 5570 3302 5582 3358
rect 5638 3302 5650 3358
rect 5570 3268 5650 3302
rect 5570 3212 5582 3268
rect 5638 3212 5650 3268
rect 5570 3178 5650 3212
rect 5570 3122 5582 3178
rect 5638 3122 5650 3178
rect 5570 3110 5650 3122
rect 5870 3628 5950 3650
rect 5870 3572 5882 3628
rect 5938 3572 5950 3628
rect 5870 3538 5950 3572
rect 5870 3482 5882 3538
rect 5938 3482 5950 3538
rect 5870 3448 5950 3482
rect 5870 3392 5882 3448
rect 5938 3392 5950 3448
rect 5870 3358 5950 3392
rect 5870 3302 5882 3358
rect 5938 3302 5950 3358
rect 5870 3268 5950 3302
rect 5870 3212 5882 3268
rect 5938 3212 5950 3268
rect 5870 3178 5950 3212
rect 5870 3122 5882 3178
rect 5938 3122 5950 3178
rect 5870 3110 5950 3122
rect 6170 3628 6250 3650
rect 6170 3572 6182 3628
rect 6238 3572 6250 3628
rect 6170 3538 6250 3572
rect 6170 3482 6182 3538
rect 6238 3482 6250 3538
rect 6170 3448 6250 3482
rect 6170 3392 6182 3448
rect 6238 3392 6250 3448
rect 6170 3358 6250 3392
rect 6170 3302 6182 3358
rect 6238 3302 6250 3358
rect 6170 3268 6250 3302
rect 6170 3212 6182 3268
rect 6238 3212 6250 3268
rect 6170 3178 6250 3212
rect 6170 3122 6182 3178
rect 6238 3122 6250 3178
rect 6170 3110 6250 3122
rect -70 2518 10 2530
rect -70 2462 -58 2518
rect -2 2462 10 2518
rect -210 2428 -130 2440
rect -210 2372 -198 2428
rect -142 2372 -130 2428
rect -210 2338 -130 2372
rect -70 2428 10 2462
rect -70 2372 -58 2428
rect -2 2420 10 2428
rect 6570 2518 6650 2530
rect 6570 2462 6582 2518
rect 6638 2462 6650 2518
rect 6570 2428 6650 2462
rect 6570 2420 6582 2428
rect -2 2416 2560 2420
rect -2 2372 1589 2416
rect -70 2364 1589 2372
rect 1641 2364 1889 2416
rect 1941 2364 2189 2416
rect 2241 2364 2489 2416
rect 2541 2364 2560 2416
rect -70 2360 2560 2364
rect 3970 2416 6582 2420
rect 3970 2364 3989 2416
rect 4041 2364 4289 2416
rect 4341 2364 4589 2416
rect 4641 2364 4889 2416
rect 4941 2372 6582 2416
rect 6638 2372 6650 2428
rect 4941 2364 6650 2372
rect 3970 2360 6650 2364
rect 6710 2428 6790 2440
rect 6710 2372 6722 2428
rect 6778 2372 6790 2428
rect -210 2282 -198 2338
rect -142 2330 -130 2338
rect 6710 2338 6790 2372
rect 6710 2330 6722 2338
rect -142 2326 1350 2330
rect -142 2282 379 2326
rect -210 2274 379 2282
rect 431 2274 679 2326
rect 731 2274 979 2326
rect 1031 2274 1279 2326
rect 1331 2274 1350 2326
rect -210 2270 1350 2274
rect 5170 2326 6722 2330
rect 5170 2274 5189 2326
rect 5241 2274 5489 2326
rect 5541 2274 5789 2326
rect 5841 2274 6089 2326
rect 6141 2282 6722 2326
rect 6778 2282 6790 2338
rect 6141 2274 6790 2282
rect 5170 2270 6790 2274
rect 1560 2236 6660 2240
rect -70 2226 10 2230
rect -70 2174 -56 2226
rect -4 2174 10 2226
rect 1560 2184 1589 2236
rect 1641 2184 1889 2236
rect 1941 2184 2189 2236
rect 2241 2184 2489 2236
rect 2541 2184 3989 2236
rect 4041 2184 4289 2236
rect 4341 2184 4589 2236
rect 4641 2184 4889 2236
rect 4941 2184 6514 2236
rect 6566 2184 6594 2236
rect 6646 2184 6660 2236
rect 1560 2180 6660 2184
rect -70 2150 10 2174
rect -70 2146 1350 2150
rect -70 2094 -56 2146
rect -4 2094 379 2146
rect 431 2094 679 2146
rect 731 2094 979 2146
rect 1031 2094 1279 2146
rect 1331 2094 1350 2146
rect -70 2090 1350 2094
rect 2770 2146 3760 2150
rect 2770 2094 2789 2146
rect 2841 2094 3089 2146
rect 3141 2094 3389 2146
rect 3441 2094 3689 2146
rect 3741 2094 3760 2146
rect 2770 2090 3760 2094
rect 5170 2146 6790 2150
rect 5170 2094 5189 2146
rect 5241 2094 5489 2146
rect 5541 2094 5789 2146
rect 5841 2094 6089 2146
rect 6141 2094 6644 2146
rect 6696 2094 6724 2146
rect 6776 2094 6790 2146
rect 5170 2090 6790 2094
rect 470 1318 550 1340
rect 470 1262 482 1318
rect 538 1262 550 1318
rect 470 1228 550 1262
rect 470 1172 482 1228
rect 538 1172 550 1228
rect 470 1138 550 1172
rect 470 1082 482 1138
rect 538 1082 550 1138
rect 470 1048 550 1082
rect 470 992 482 1048
rect 538 992 550 1048
rect 470 958 550 992
rect 470 902 482 958
rect 538 902 550 958
rect 470 868 550 902
rect 470 812 482 868
rect 538 812 550 868
rect 470 800 550 812
rect 770 1318 850 1340
rect 770 1262 782 1318
rect 838 1262 850 1318
rect 770 1228 850 1262
rect 770 1172 782 1228
rect 838 1172 850 1228
rect 770 1138 850 1172
rect 770 1082 782 1138
rect 838 1082 850 1138
rect 770 1048 850 1082
rect 770 992 782 1048
rect 838 992 850 1048
rect 770 958 850 992
rect 770 902 782 958
rect 838 902 850 958
rect 770 868 850 902
rect 770 812 782 868
rect 838 812 850 868
rect 770 800 850 812
rect 1070 1318 1150 1340
rect 1070 1262 1082 1318
rect 1138 1262 1150 1318
rect 1070 1228 1150 1262
rect 1070 1172 1082 1228
rect 1138 1172 1150 1228
rect 1070 1138 1150 1172
rect 1070 1082 1082 1138
rect 1138 1082 1150 1138
rect 1070 1048 1150 1082
rect 1070 992 1082 1048
rect 1138 992 1150 1048
rect 1070 958 1150 992
rect 1070 902 1082 958
rect 1138 902 1150 958
rect 1070 868 1150 902
rect 1070 812 1082 868
rect 1138 812 1150 868
rect 1070 800 1150 812
rect 1370 1318 1450 1340
rect 1370 1262 1382 1318
rect 1438 1262 1450 1318
rect 1370 1228 1450 1262
rect 1370 1172 1382 1228
rect 1438 1172 1450 1228
rect 1370 1138 1450 1172
rect 1370 1082 1382 1138
rect 1438 1082 1450 1138
rect 1370 1048 1450 1082
rect 1370 992 1382 1048
rect 1438 992 1450 1048
rect 1370 958 1450 992
rect 1370 902 1382 958
rect 1438 902 1450 958
rect 1370 868 1450 902
rect 1370 812 1382 868
rect 1438 812 1450 868
rect 1370 800 1450 812
rect 1670 1318 1750 1340
rect 1670 1262 1682 1318
rect 1738 1262 1750 1318
rect 1670 1228 1750 1262
rect 1670 1172 1682 1228
rect 1738 1172 1750 1228
rect 1670 1138 1750 1172
rect 1670 1082 1682 1138
rect 1738 1082 1750 1138
rect 1670 1048 1750 1082
rect 1670 992 1682 1048
rect 1738 992 1750 1048
rect 1670 958 1750 992
rect 1670 902 1682 958
rect 1738 902 1750 958
rect 1670 868 1750 902
rect 1670 812 1682 868
rect 1738 812 1750 868
rect 1670 800 1750 812
rect 1970 1318 2050 1340
rect 1970 1262 1982 1318
rect 2038 1262 2050 1318
rect 1970 1228 2050 1262
rect 1970 1172 1982 1228
rect 2038 1172 2050 1228
rect 1970 1138 2050 1172
rect 1970 1082 1982 1138
rect 2038 1082 2050 1138
rect 1970 1048 2050 1082
rect 1970 992 1982 1048
rect 2038 992 2050 1048
rect 1970 958 2050 992
rect 1970 902 1982 958
rect 2038 902 2050 958
rect 1970 868 2050 902
rect 1970 812 1982 868
rect 2038 812 2050 868
rect 1970 800 2050 812
rect 2270 1318 2350 1340
rect 2270 1262 2282 1318
rect 2338 1262 2350 1318
rect 2270 1228 2350 1262
rect 2270 1172 2282 1228
rect 2338 1172 2350 1228
rect 2270 1138 2350 1172
rect 2270 1082 2282 1138
rect 2338 1082 2350 1138
rect 2270 1048 2350 1082
rect 2270 992 2282 1048
rect 2338 992 2350 1048
rect 2270 958 2350 992
rect 2270 902 2282 958
rect 2338 902 2350 958
rect 2270 868 2350 902
rect 2270 812 2282 868
rect 2338 812 2350 868
rect 2270 800 2350 812
rect 2570 1318 2650 1340
rect 2570 1262 2582 1318
rect 2638 1262 2650 1318
rect 2570 1228 2650 1262
rect 2570 1172 2582 1228
rect 2638 1172 2650 1228
rect 2570 1138 2650 1172
rect 2570 1082 2582 1138
rect 2638 1082 2650 1138
rect 2570 1048 2650 1082
rect 2570 992 2582 1048
rect 2638 992 2650 1048
rect 2570 958 2650 992
rect 2570 902 2582 958
rect 2638 902 2650 958
rect 2570 868 2650 902
rect 2570 812 2582 868
rect 2638 812 2650 868
rect 2570 800 2650 812
rect 2870 1318 2950 1340
rect 2870 1262 2882 1318
rect 2938 1262 2950 1318
rect 2870 1228 2950 1262
rect 2870 1172 2882 1228
rect 2938 1172 2950 1228
rect 2870 1138 2950 1172
rect 2870 1082 2882 1138
rect 2938 1082 2950 1138
rect 2870 1048 2950 1082
rect 2870 992 2882 1048
rect 2938 992 2950 1048
rect 2870 958 2950 992
rect 2870 902 2882 958
rect 2938 902 2950 958
rect 2870 868 2950 902
rect 2870 812 2882 868
rect 2938 812 2950 868
rect 2870 800 2950 812
rect 3470 1318 3550 1340
rect 3470 1262 3482 1318
rect 3538 1262 3550 1318
rect 3470 1228 3550 1262
rect 3470 1172 3482 1228
rect 3538 1172 3550 1228
rect 3470 1138 3550 1172
rect 3470 1082 3482 1138
rect 3538 1082 3550 1138
rect 3470 1048 3550 1082
rect 3470 992 3482 1048
rect 3538 992 3550 1048
rect 3470 958 3550 992
rect 3470 902 3482 958
rect 3538 902 3550 958
rect 3470 868 3550 902
rect 3470 812 3482 868
rect 3538 812 3550 868
rect 3470 800 3550 812
rect 3770 1318 3850 1340
rect 3770 1262 3782 1318
rect 3838 1262 3850 1318
rect 3770 1228 3850 1262
rect 3770 1172 3782 1228
rect 3838 1172 3850 1228
rect 3770 1138 3850 1172
rect 3770 1082 3782 1138
rect 3838 1082 3850 1138
rect 3770 1048 3850 1082
rect 3770 992 3782 1048
rect 3838 992 3850 1048
rect 3770 958 3850 992
rect 3770 902 3782 958
rect 3838 902 3850 958
rect 3770 868 3850 902
rect 3770 812 3782 868
rect 3838 812 3850 868
rect 3770 800 3850 812
rect 4070 1318 4150 1340
rect 4070 1262 4082 1318
rect 4138 1262 4150 1318
rect 4070 1228 4150 1262
rect 4070 1172 4082 1228
rect 4138 1172 4150 1228
rect 4070 1138 4150 1172
rect 4070 1082 4082 1138
rect 4138 1082 4150 1138
rect 4070 1048 4150 1082
rect 4070 992 4082 1048
rect 4138 992 4150 1048
rect 4070 958 4150 992
rect 4070 902 4082 958
rect 4138 902 4150 958
rect 4070 868 4150 902
rect 4070 812 4082 868
rect 4138 812 4150 868
rect 4070 800 4150 812
rect 4370 1318 4450 1340
rect 4370 1262 4382 1318
rect 4438 1262 4450 1318
rect 4370 1228 4450 1262
rect 4370 1172 4382 1228
rect 4438 1172 4450 1228
rect 4370 1138 4450 1172
rect 4370 1082 4382 1138
rect 4438 1082 4450 1138
rect 4370 1048 4450 1082
rect 4370 992 4382 1048
rect 4438 992 4450 1048
rect 4370 958 4450 992
rect 4370 902 4382 958
rect 4438 902 4450 958
rect 4370 868 4450 902
rect 4370 812 4382 868
rect 4438 812 4450 868
rect 4370 800 4450 812
rect 4670 1318 4750 1340
rect 4670 1262 4682 1318
rect 4738 1262 4750 1318
rect 4670 1228 4750 1262
rect 4670 1172 4682 1228
rect 4738 1172 4750 1228
rect 4670 1138 4750 1172
rect 4670 1082 4682 1138
rect 4738 1082 4750 1138
rect 4670 1048 4750 1082
rect 4670 992 4682 1048
rect 4738 992 4750 1048
rect 4670 958 4750 992
rect 4670 902 4682 958
rect 4738 902 4750 958
rect 4670 868 4750 902
rect 4670 812 4682 868
rect 4738 812 4750 868
rect 4670 800 4750 812
rect 4970 1318 5050 1340
rect 4970 1262 4982 1318
rect 5038 1262 5050 1318
rect 4970 1228 5050 1262
rect 4970 1172 4982 1228
rect 5038 1172 5050 1228
rect 4970 1138 5050 1172
rect 4970 1082 4982 1138
rect 5038 1082 5050 1138
rect 4970 1048 5050 1082
rect 4970 992 4982 1048
rect 5038 992 5050 1048
rect 4970 958 5050 992
rect 4970 902 4982 958
rect 5038 902 5050 958
rect 4970 868 5050 902
rect 4970 812 4982 868
rect 5038 812 5050 868
rect 4970 800 5050 812
rect 5270 1318 5350 1340
rect 5270 1262 5282 1318
rect 5338 1262 5350 1318
rect 5270 1228 5350 1262
rect 5270 1172 5282 1228
rect 5338 1172 5350 1228
rect 5270 1138 5350 1172
rect 5270 1082 5282 1138
rect 5338 1082 5350 1138
rect 5270 1048 5350 1082
rect 5270 992 5282 1048
rect 5338 992 5350 1048
rect 5270 958 5350 992
rect 5270 902 5282 958
rect 5338 902 5350 958
rect 5270 868 5350 902
rect 5270 812 5282 868
rect 5338 812 5350 868
rect 5270 800 5350 812
rect 5570 1318 5650 1340
rect 5570 1262 5582 1318
rect 5638 1262 5650 1318
rect 5570 1228 5650 1262
rect 5570 1172 5582 1228
rect 5638 1172 5650 1228
rect 5570 1138 5650 1172
rect 5570 1082 5582 1138
rect 5638 1082 5650 1138
rect 5570 1048 5650 1082
rect 5570 992 5582 1048
rect 5638 992 5650 1048
rect 5570 958 5650 992
rect 5570 902 5582 958
rect 5638 902 5650 958
rect 5570 868 5650 902
rect 5570 812 5582 868
rect 5638 812 5650 868
rect 5570 800 5650 812
rect 5870 1318 5950 1340
rect 5870 1262 5882 1318
rect 5938 1262 5950 1318
rect 5870 1228 5950 1262
rect 5870 1172 5882 1228
rect 5938 1172 5950 1228
rect 5870 1138 5950 1172
rect 5870 1082 5882 1138
rect 5938 1082 5950 1138
rect 5870 1048 5950 1082
rect 5870 992 5882 1048
rect 5938 992 5950 1048
rect 5870 958 5950 992
rect 5870 902 5882 958
rect 5938 902 5950 958
rect 5870 868 5950 902
rect 5870 812 5882 868
rect 5938 812 5950 868
rect 5870 800 5950 812
rect 6170 1318 6250 1340
rect 6170 1262 6182 1318
rect 6238 1262 6250 1318
rect 6170 1228 6250 1262
rect 6170 1172 6182 1228
rect 6238 1172 6250 1228
rect 6170 1138 6250 1172
rect 6170 1082 6182 1138
rect 6238 1082 6250 1138
rect 6170 1048 6250 1082
rect 6170 992 6182 1048
rect 6238 992 6250 1048
rect 6170 958 6250 992
rect 6170 902 6182 958
rect 6238 902 6250 958
rect 6170 868 6250 902
rect 6170 812 6182 868
rect 6238 812 6250 868
rect 6170 800 6250 812
rect -70 198 10 210
rect -70 142 -58 198
rect -2 142 10 198
rect -210 108 -130 120
rect -210 52 -198 108
rect -142 52 -130 108
rect -210 18 -130 52
rect -70 108 10 142
rect -70 52 -58 108
rect -2 100 10 108
rect 6570 198 6650 210
rect 6570 142 6582 198
rect 6638 142 6650 198
rect 6570 108 6650 142
rect 6570 100 6582 108
rect -2 96 1350 100
rect -2 52 379 96
rect -70 44 379 52
rect 431 44 679 96
rect 731 44 979 96
rect 1031 44 1279 96
rect 1331 44 1350 96
rect -70 40 1350 44
rect 5170 96 6582 100
rect 5170 44 5189 96
rect 5241 44 5489 96
rect 5541 44 5789 96
rect 5841 44 6089 96
rect 6141 52 6582 96
rect 6638 52 6650 108
rect 6141 44 6650 52
rect 5170 40 6650 44
rect 6710 108 6790 120
rect 6710 52 6722 108
rect 6778 52 6790 108
rect -210 -38 -198 18
rect -142 10 -130 18
rect 6710 18 6790 52
rect 6710 10 6722 18
rect -142 6 2550 10
rect -142 -38 1579 6
rect -210 -46 1579 -38
rect 1631 -46 1879 6
rect 1931 -46 2179 6
rect 2231 -46 2479 6
rect 2531 -46 2550 6
rect -210 -50 2550 -46
rect 3970 6 6722 10
rect 3970 -46 3989 6
rect 4041 -46 4289 6
rect 4341 -46 4589 6
rect 4641 -46 4889 6
rect 4941 -38 6722 6
rect 6778 -38 6790 18
rect 4941 -46 6790 -38
rect 3970 -50 6790 -46
rect -70 -222 10 -210
rect -70 -278 -58 -222
rect -2 -278 10 -222
rect -210 -312 -130 -300
rect -210 -368 -198 -312
rect -142 -368 -130 -312
rect -210 -402 -130 -368
rect -70 -312 10 -278
rect -70 -368 -58 -312
rect -2 -320 10 -312
rect 6570 -222 6650 -210
rect 6570 -278 6582 -222
rect 6638 -278 6650 -222
rect 6570 -312 6650 -278
rect 6570 -320 6582 -312
rect -2 -368 6582 -320
rect 6638 -368 6650 -312
rect -70 -380 6650 -368
rect 6710 -312 6790 -300
rect 6710 -368 6722 -312
rect 6778 -368 6790 -312
rect -210 -458 -198 -402
rect -142 -410 -130 -402
rect 6710 -402 6790 -368
rect 6710 -410 6722 -402
rect -142 -458 6722 -410
rect 6778 -458 6790 -402
rect -210 -470 6790 -458
<< via2 >>
rect 6494 5266 6550 5268
rect 6494 5214 6496 5266
rect 6496 5214 6548 5266
rect 6548 5214 6550 5266
rect 6494 5212 6550 5214
rect 6734 5212 6790 5268
rect 482 3626 538 3628
rect 482 3574 484 3626
rect 484 3574 536 3626
rect 536 3574 538 3626
rect 482 3572 538 3574
rect 482 3536 538 3538
rect 482 3484 484 3536
rect 484 3484 536 3536
rect 536 3484 538 3536
rect 482 3482 538 3484
rect 482 3446 538 3448
rect 482 3394 484 3446
rect 484 3394 536 3446
rect 536 3394 538 3446
rect 482 3392 538 3394
rect 482 3356 538 3358
rect 482 3304 484 3356
rect 484 3304 536 3356
rect 536 3304 538 3356
rect 482 3302 538 3304
rect 482 3266 538 3268
rect 482 3214 484 3266
rect 484 3214 536 3266
rect 536 3214 538 3266
rect 482 3212 538 3214
rect 482 3176 538 3178
rect 482 3124 484 3176
rect 484 3124 536 3176
rect 536 3124 538 3176
rect 482 3122 538 3124
rect 782 3626 838 3628
rect 782 3574 784 3626
rect 784 3574 836 3626
rect 836 3574 838 3626
rect 782 3572 838 3574
rect 782 3536 838 3538
rect 782 3484 784 3536
rect 784 3484 836 3536
rect 836 3484 838 3536
rect 782 3482 838 3484
rect 782 3446 838 3448
rect 782 3394 784 3446
rect 784 3394 836 3446
rect 836 3394 838 3446
rect 782 3392 838 3394
rect 782 3356 838 3358
rect 782 3304 784 3356
rect 784 3304 836 3356
rect 836 3304 838 3356
rect 782 3302 838 3304
rect 782 3266 838 3268
rect 782 3214 784 3266
rect 784 3214 836 3266
rect 836 3214 838 3266
rect 782 3212 838 3214
rect 782 3176 838 3178
rect 782 3124 784 3176
rect 784 3124 836 3176
rect 836 3124 838 3176
rect 782 3122 838 3124
rect 1082 3626 1138 3628
rect 1082 3574 1084 3626
rect 1084 3574 1136 3626
rect 1136 3574 1138 3626
rect 1082 3572 1138 3574
rect 1082 3536 1138 3538
rect 1082 3484 1084 3536
rect 1084 3484 1136 3536
rect 1136 3484 1138 3536
rect 1082 3482 1138 3484
rect 1082 3446 1138 3448
rect 1082 3394 1084 3446
rect 1084 3394 1136 3446
rect 1136 3394 1138 3446
rect 1082 3392 1138 3394
rect 1082 3356 1138 3358
rect 1082 3304 1084 3356
rect 1084 3304 1136 3356
rect 1136 3304 1138 3356
rect 1082 3302 1138 3304
rect 1082 3266 1138 3268
rect 1082 3214 1084 3266
rect 1084 3214 1136 3266
rect 1136 3214 1138 3266
rect 1082 3212 1138 3214
rect 1082 3176 1138 3178
rect 1082 3124 1084 3176
rect 1084 3124 1136 3176
rect 1136 3124 1138 3176
rect 1082 3122 1138 3124
rect 1382 3626 1438 3628
rect 1382 3574 1384 3626
rect 1384 3574 1436 3626
rect 1436 3574 1438 3626
rect 1382 3572 1438 3574
rect 1382 3536 1438 3538
rect 1382 3484 1384 3536
rect 1384 3484 1436 3536
rect 1436 3484 1438 3536
rect 1382 3482 1438 3484
rect 1382 3446 1438 3448
rect 1382 3394 1384 3446
rect 1384 3394 1436 3446
rect 1436 3394 1438 3446
rect 1382 3392 1438 3394
rect 1382 3356 1438 3358
rect 1382 3304 1384 3356
rect 1384 3304 1436 3356
rect 1436 3304 1438 3356
rect 1382 3302 1438 3304
rect 1382 3266 1438 3268
rect 1382 3214 1384 3266
rect 1384 3214 1436 3266
rect 1436 3214 1438 3266
rect 1382 3212 1438 3214
rect 1382 3176 1438 3178
rect 1382 3124 1384 3176
rect 1384 3124 1436 3176
rect 1436 3124 1438 3176
rect 1382 3122 1438 3124
rect 1682 3626 1738 3628
rect 1682 3574 1684 3626
rect 1684 3574 1736 3626
rect 1736 3574 1738 3626
rect 1682 3572 1738 3574
rect 1682 3536 1738 3538
rect 1682 3484 1684 3536
rect 1684 3484 1736 3536
rect 1736 3484 1738 3536
rect 1682 3482 1738 3484
rect 1682 3446 1738 3448
rect 1682 3394 1684 3446
rect 1684 3394 1736 3446
rect 1736 3394 1738 3446
rect 1682 3392 1738 3394
rect 1682 3356 1738 3358
rect 1682 3304 1684 3356
rect 1684 3304 1736 3356
rect 1736 3304 1738 3356
rect 1682 3302 1738 3304
rect 1682 3266 1738 3268
rect 1682 3214 1684 3266
rect 1684 3214 1736 3266
rect 1736 3214 1738 3266
rect 1682 3212 1738 3214
rect 1682 3176 1738 3178
rect 1682 3124 1684 3176
rect 1684 3124 1736 3176
rect 1736 3124 1738 3176
rect 1682 3122 1738 3124
rect 1982 3626 2038 3628
rect 1982 3574 1984 3626
rect 1984 3574 2036 3626
rect 2036 3574 2038 3626
rect 1982 3572 2038 3574
rect 1982 3536 2038 3538
rect 1982 3484 1984 3536
rect 1984 3484 2036 3536
rect 2036 3484 2038 3536
rect 1982 3482 2038 3484
rect 1982 3446 2038 3448
rect 1982 3394 1984 3446
rect 1984 3394 2036 3446
rect 2036 3394 2038 3446
rect 1982 3392 2038 3394
rect 1982 3356 2038 3358
rect 1982 3304 1984 3356
rect 1984 3304 2036 3356
rect 2036 3304 2038 3356
rect 1982 3302 2038 3304
rect 1982 3266 2038 3268
rect 1982 3214 1984 3266
rect 1984 3214 2036 3266
rect 2036 3214 2038 3266
rect 1982 3212 2038 3214
rect 1982 3176 2038 3178
rect 1982 3124 1984 3176
rect 1984 3124 2036 3176
rect 2036 3124 2038 3176
rect 1982 3122 2038 3124
rect 2282 3626 2338 3628
rect 2282 3574 2284 3626
rect 2284 3574 2336 3626
rect 2336 3574 2338 3626
rect 2282 3572 2338 3574
rect 2282 3536 2338 3538
rect 2282 3484 2284 3536
rect 2284 3484 2336 3536
rect 2336 3484 2338 3536
rect 2282 3482 2338 3484
rect 2282 3446 2338 3448
rect 2282 3394 2284 3446
rect 2284 3394 2336 3446
rect 2336 3394 2338 3446
rect 2282 3392 2338 3394
rect 2282 3356 2338 3358
rect 2282 3304 2284 3356
rect 2284 3304 2336 3356
rect 2336 3304 2338 3356
rect 2282 3302 2338 3304
rect 2282 3266 2338 3268
rect 2282 3214 2284 3266
rect 2284 3214 2336 3266
rect 2336 3214 2338 3266
rect 2282 3212 2338 3214
rect 2282 3176 2338 3178
rect 2282 3124 2284 3176
rect 2284 3124 2336 3176
rect 2336 3124 2338 3176
rect 2282 3122 2338 3124
rect 2582 3626 2638 3628
rect 2582 3574 2584 3626
rect 2584 3574 2636 3626
rect 2636 3574 2638 3626
rect 2582 3572 2638 3574
rect 2582 3536 2638 3538
rect 2582 3484 2584 3536
rect 2584 3484 2636 3536
rect 2636 3484 2638 3536
rect 2582 3482 2638 3484
rect 2582 3446 2638 3448
rect 2582 3394 2584 3446
rect 2584 3394 2636 3446
rect 2636 3394 2638 3446
rect 2582 3392 2638 3394
rect 2582 3356 2638 3358
rect 2582 3304 2584 3356
rect 2584 3304 2636 3356
rect 2636 3304 2638 3356
rect 2582 3302 2638 3304
rect 2582 3266 2638 3268
rect 2582 3214 2584 3266
rect 2584 3214 2636 3266
rect 2636 3214 2638 3266
rect 2582 3212 2638 3214
rect 2582 3176 2638 3178
rect 2582 3124 2584 3176
rect 2584 3124 2636 3176
rect 2636 3124 2638 3176
rect 2582 3122 2638 3124
rect 2882 3626 2938 3628
rect 2882 3574 2884 3626
rect 2884 3574 2936 3626
rect 2936 3574 2938 3626
rect 2882 3572 2938 3574
rect 2882 3536 2938 3538
rect 2882 3484 2884 3536
rect 2884 3484 2936 3536
rect 2936 3484 2938 3536
rect 2882 3482 2938 3484
rect 2882 3446 2938 3448
rect 2882 3394 2884 3446
rect 2884 3394 2936 3446
rect 2936 3394 2938 3446
rect 2882 3392 2938 3394
rect 2882 3356 2938 3358
rect 2882 3304 2884 3356
rect 2884 3304 2936 3356
rect 2936 3304 2938 3356
rect 2882 3302 2938 3304
rect 2882 3266 2938 3268
rect 2882 3214 2884 3266
rect 2884 3214 2936 3266
rect 2936 3214 2938 3266
rect 2882 3212 2938 3214
rect 2882 3176 2938 3178
rect 2882 3124 2884 3176
rect 2884 3124 2936 3176
rect 2936 3124 2938 3176
rect 2882 3122 2938 3124
rect 3182 3626 3238 3628
rect 3182 3574 3184 3626
rect 3184 3574 3236 3626
rect 3236 3574 3238 3626
rect 3182 3572 3238 3574
rect 3182 3536 3238 3538
rect 3182 3484 3184 3536
rect 3184 3484 3236 3536
rect 3236 3484 3238 3536
rect 3182 3482 3238 3484
rect 3182 3446 3238 3448
rect 3182 3394 3184 3446
rect 3184 3394 3236 3446
rect 3236 3394 3238 3446
rect 3182 3392 3238 3394
rect 3182 3356 3238 3358
rect 3182 3304 3184 3356
rect 3184 3304 3236 3356
rect 3236 3304 3238 3356
rect 3182 3302 3238 3304
rect 3182 3266 3238 3268
rect 3182 3214 3184 3266
rect 3184 3214 3236 3266
rect 3236 3214 3238 3266
rect 3182 3212 3238 3214
rect 3182 3176 3238 3178
rect 3182 3124 3184 3176
rect 3184 3124 3236 3176
rect 3236 3124 3238 3176
rect 3182 3122 3238 3124
rect 3782 3626 3838 3628
rect 3782 3574 3784 3626
rect 3784 3574 3836 3626
rect 3836 3574 3838 3626
rect 3782 3572 3838 3574
rect 3782 3536 3838 3538
rect 3782 3484 3784 3536
rect 3784 3484 3836 3536
rect 3836 3484 3838 3536
rect 3782 3482 3838 3484
rect 3782 3446 3838 3448
rect 3782 3394 3784 3446
rect 3784 3394 3836 3446
rect 3836 3394 3838 3446
rect 3782 3392 3838 3394
rect 3782 3356 3838 3358
rect 3782 3304 3784 3356
rect 3784 3304 3836 3356
rect 3836 3304 3838 3356
rect 3782 3302 3838 3304
rect 3782 3266 3838 3268
rect 3782 3214 3784 3266
rect 3784 3214 3836 3266
rect 3836 3214 3838 3266
rect 3782 3212 3838 3214
rect 3782 3176 3838 3178
rect 3782 3124 3784 3176
rect 3784 3124 3836 3176
rect 3836 3124 3838 3176
rect 3782 3122 3838 3124
rect 4082 3626 4138 3628
rect 4082 3574 4084 3626
rect 4084 3574 4136 3626
rect 4136 3574 4138 3626
rect 4082 3572 4138 3574
rect 4082 3536 4138 3538
rect 4082 3484 4084 3536
rect 4084 3484 4136 3536
rect 4136 3484 4138 3536
rect 4082 3482 4138 3484
rect 4082 3446 4138 3448
rect 4082 3394 4084 3446
rect 4084 3394 4136 3446
rect 4136 3394 4138 3446
rect 4082 3392 4138 3394
rect 4082 3356 4138 3358
rect 4082 3304 4084 3356
rect 4084 3304 4136 3356
rect 4136 3304 4138 3356
rect 4082 3302 4138 3304
rect 4082 3266 4138 3268
rect 4082 3214 4084 3266
rect 4084 3214 4136 3266
rect 4136 3214 4138 3266
rect 4082 3212 4138 3214
rect 4082 3176 4138 3178
rect 4082 3124 4084 3176
rect 4084 3124 4136 3176
rect 4136 3124 4138 3176
rect 4082 3122 4138 3124
rect 4382 3626 4438 3628
rect 4382 3574 4384 3626
rect 4384 3574 4436 3626
rect 4436 3574 4438 3626
rect 4382 3572 4438 3574
rect 4382 3536 4438 3538
rect 4382 3484 4384 3536
rect 4384 3484 4436 3536
rect 4436 3484 4438 3536
rect 4382 3482 4438 3484
rect 4382 3446 4438 3448
rect 4382 3394 4384 3446
rect 4384 3394 4436 3446
rect 4436 3394 4438 3446
rect 4382 3392 4438 3394
rect 4382 3356 4438 3358
rect 4382 3304 4384 3356
rect 4384 3304 4436 3356
rect 4436 3304 4438 3356
rect 4382 3302 4438 3304
rect 4382 3266 4438 3268
rect 4382 3214 4384 3266
rect 4384 3214 4436 3266
rect 4436 3214 4438 3266
rect 4382 3212 4438 3214
rect 4382 3176 4438 3178
rect 4382 3124 4384 3176
rect 4384 3124 4436 3176
rect 4436 3124 4438 3176
rect 4382 3122 4438 3124
rect 4682 3626 4738 3628
rect 4682 3574 4684 3626
rect 4684 3574 4736 3626
rect 4736 3574 4738 3626
rect 4682 3572 4738 3574
rect 4682 3536 4738 3538
rect 4682 3484 4684 3536
rect 4684 3484 4736 3536
rect 4736 3484 4738 3536
rect 4682 3482 4738 3484
rect 4682 3446 4738 3448
rect 4682 3394 4684 3446
rect 4684 3394 4736 3446
rect 4736 3394 4738 3446
rect 4682 3392 4738 3394
rect 4682 3356 4738 3358
rect 4682 3304 4684 3356
rect 4684 3304 4736 3356
rect 4736 3304 4738 3356
rect 4682 3302 4738 3304
rect 4682 3266 4738 3268
rect 4682 3214 4684 3266
rect 4684 3214 4736 3266
rect 4736 3214 4738 3266
rect 4682 3212 4738 3214
rect 4682 3176 4738 3178
rect 4682 3124 4684 3176
rect 4684 3124 4736 3176
rect 4736 3124 4738 3176
rect 4682 3122 4738 3124
rect 4982 3626 5038 3628
rect 4982 3574 4984 3626
rect 4984 3574 5036 3626
rect 5036 3574 5038 3626
rect 4982 3572 5038 3574
rect 4982 3536 5038 3538
rect 4982 3484 4984 3536
rect 4984 3484 5036 3536
rect 5036 3484 5038 3536
rect 4982 3482 5038 3484
rect 4982 3446 5038 3448
rect 4982 3394 4984 3446
rect 4984 3394 5036 3446
rect 5036 3394 5038 3446
rect 4982 3392 5038 3394
rect 4982 3356 5038 3358
rect 4982 3304 4984 3356
rect 4984 3304 5036 3356
rect 5036 3304 5038 3356
rect 4982 3302 5038 3304
rect 4982 3266 5038 3268
rect 4982 3214 4984 3266
rect 4984 3214 5036 3266
rect 5036 3214 5038 3266
rect 4982 3212 5038 3214
rect 4982 3176 5038 3178
rect 4982 3124 4984 3176
rect 4984 3124 5036 3176
rect 5036 3124 5038 3176
rect 4982 3122 5038 3124
rect 5282 3626 5338 3628
rect 5282 3574 5284 3626
rect 5284 3574 5336 3626
rect 5336 3574 5338 3626
rect 5282 3572 5338 3574
rect 5282 3536 5338 3538
rect 5282 3484 5284 3536
rect 5284 3484 5336 3536
rect 5336 3484 5338 3536
rect 5282 3482 5338 3484
rect 5282 3446 5338 3448
rect 5282 3394 5284 3446
rect 5284 3394 5336 3446
rect 5336 3394 5338 3446
rect 5282 3392 5338 3394
rect 5282 3356 5338 3358
rect 5282 3304 5284 3356
rect 5284 3304 5336 3356
rect 5336 3304 5338 3356
rect 5282 3302 5338 3304
rect 5282 3266 5338 3268
rect 5282 3214 5284 3266
rect 5284 3214 5336 3266
rect 5336 3214 5338 3266
rect 5282 3212 5338 3214
rect 5282 3176 5338 3178
rect 5282 3124 5284 3176
rect 5284 3124 5336 3176
rect 5336 3124 5338 3176
rect 5282 3122 5338 3124
rect 5582 3626 5638 3628
rect 5582 3574 5584 3626
rect 5584 3574 5636 3626
rect 5636 3574 5638 3626
rect 5582 3572 5638 3574
rect 5582 3536 5638 3538
rect 5582 3484 5584 3536
rect 5584 3484 5636 3536
rect 5636 3484 5638 3536
rect 5582 3482 5638 3484
rect 5582 3446 5638 3448
rect 5582 3394 5584 3446
rect 5584 3394 5636 3446
rect 5636 3394 5638 3446
rect 5582 3392 5638 3394
rect 5582 3356 5638 3358
rect 5582 3304 5584 3356
rect 5584 3304 5636 3356
rect 5636 3304 5638 3356
rect 5582 3302 5638 3304
rect 5582 3266 5638 3268
rect 5582 3214 5584 3266
rect 5584 3214 5636 3266
rect 5636 3214 5638 3266
rect 5582 3212 5638 3214
rect 5582 3176 5638 3178
rect 5582 3124 5584 3176
rect 5584 3124 5636 3176
rect 5636 3124 5638 3176
rect 5582 3122 5638 3124
rect 5882 3626 5938 3628
rect 5882 3574 5884 3626
rect 5884 3574 5936 3626
rect 5936 3574 5938 3626
rect 5882 3572 5938 3574
rect 5882 3536 5938 3538
rect 5882 3484 5884 3536
rect 5884 3484 5936 3536
rect 5936 3484 5938 3536
rect 5882 3482 5938 3484
rect 5882 3446 5938 3448
rect 5882 3394 5884 3446
rect 5884 3394 5936 3446
rect 5936 3394 5938 3446
rect 5882 3392 5938 3394
rect 5882 3356 5938 3358
rect 5882 3304 5884 3356
rect 5884 3304 5936 3356
rect 5936 3304 5938 3356
rect 5882 3302 5938 3304
rect 5882 3266 5938 3268
rect 5882 3214 5884 3266
rect 5884 3214 5936 3266
rect 5936 3214 5938 3266
rect 5882 3212 5938 3214
rect 5882 3176 5938 3178
rect 5882 3124 5884 3176
rect 5884 3124 5936 3176
rect 5936 3124 5938 3176
rect 5882 3122 5938 3124
rect 6182 3626 6238 3628
rect 6182 3574 6184 3626
rect 6184 3574 6236 3626
rect 6236 3574 6238 3626
rect 6182 3572 6238 3574
rect 6182 3536 6238 3538
rect 6182 3484 6184 3536
rect 6184 3484 6236 3536
rect 6236 3484 6238 3536
rect 6182 3482 6238 3484
rect 6182 3446 6238 3448
rect 6182 3394 6184 3446
rect 6184 3394 6236 3446
rect 6236 3394 6238 3446
rect 6182 3392 6238 3394
rect 6182 3356 6238 3358
rect 6182 3304 6184 3356
rect 6184 3304 6236 3356
rect 6236 3304 6238 3356
rect 6182 3302 6238 3304
rect 6182 3266 6238 3268
rect 6182 3214 6184 3266
rect 6184 3214 6236 3266
rect 6236 3214 6238 3266
rect 6182 3212 6238 3214
rect 6182 3176 6238 3178
rect 6182 3124 6184 3176
rect 6184 3124 6236 3176
rect 6236 3124 6238 3176
rect 6182 3122 6238 3124
rect -58 2462 -2 2518
rect -198 2372 -142 2428
rect -58 2372 -2 2428
rect 6582 2462 6638 2518
rect 6582 2372 6638 2428
rect 6722 2372 6778 2428
rect -198 2282 -142 2338
rect 6722 2282 6778 2338
rect 482 1316 538 1318
rect 482 1264 484 1316
rect 484 1264 536 1316
rect 536 1264 538 1316
rect 482 1262 538 1264
rect 482 1226 538 1228
rect 482 1174 484 1226
rect 484 1174 536 1226
rect 536 1174 538 1226
rect 482 1172 538 1174
rect 482 1136 538 1138
rect 482 1084 484 1136
rect 484 1084 536 1136
rect 536 1084 538 1136
rect 482 1082 538 1084
rect 482 1046 538 1048
rect 482 994 484 1046
rect 484 994 536 1046
rect 536 994 538 1046
rect 482 992 538 994
rect 482 956 538 958
rect 482 904 484 956
rect 484 904 536 956
rect 536 904 538 956
rect 482 902 538 904
rect 482 866 538 868
rect 482 814 484 866
rect 484 814 536 866
rect 536 814 538 866
rect 482 812 538 814
rect 782 1316 838 1318
rect 782 1264 784 1316
rect 784 1264 836 1316
rect 836 1264 838 1316
rect 782 1262 838 1264
rect 782 1226 838 1228
rect 782 1174 784 1226
rect 784 1174 836 1226
rect 836 1174 838 1226
rect 782 1172 838 1174
rect 782 1136 838 1138
rect 782 1084 784 1136
rect 784 1084 836 1136
rect 836 1084 838 1136
rect 782 1082 838 1084
rect 782 1046 838 1048
rect 782 994 784 1046
rect 784 994 836 1046
rect 836 994 838 1046
rect 782 992 838 994
rect 782 956 838 958
rect 782 904 784 956
rect 784 904 836 956
rect 836 904 838 956
rect 782 902 838 904
rect 782 866 838 868
rect 782 814 784 866
rect 784 814 836 866
rect 836 814 838 866
rect 782 812 838 814
rect 1082 1316 1138 1318
rect 1082 1264 1084 1316
rect 1084 1264 1136 1316
rect 1136 1264 1138 1316
rect 1082 1262 1138 1264
rect 1082 1226 1138 1228
rect 1082 1174 1084 1226
rect 1084 1174 1136 1226
rect 1136 1174 1138 1226
rect 1082 1172 1138 1174
rect 1082 1136 1138 1138
rect 1082 1084 1084 1136
rect 1084 1084 1136 1136
rect 1136 1084 1138 1136
rect 1082 1082 1138 1084
rect 1082 1046 1138 1048
rect 1082 994 1084 1046
rect 1084 994 1136 1046
rect 1136 994 1138 1046
rect 1082 992 1138 994
rect 1082 956 1138 958
rect 1082 904 1084 956
rect 1084 904 1136 956
rect 1136 904 1138 956
rect 1082 902 1138 904
rect 1082 866 1138 868
rect 1082 814 1084 866
rect 1084 814 1136 866
rect 1136 814 1138 866
rect 1082 812 1138 814
rect 1382 1316 1438 1318
rect 1382 1264 1384 1316
rect 1384 1264 1436 1316
rect 1436 1264 1438 1316
rect 1382 1262 1438 1264
rect 1382 1226 1438 1228
rect 1382 1174 1384 1226
rect 1384 1174 1436 1226
rect 1436 1174 1438 1226
rect 1382 1172 1438 1174
rect 1382 1136 1438 1138
rect 1382 1084 1384 1136
rect 1384 1084 1436 1136
rect 1436 1084 1438 1136
rect 1382 1082 1438 1084
rect 1382 1046 1438 1048
rect 1382 994 1384 1046
rect 1384 994 1436 1046
rect 1436 994 1438 1046
rect 1382 992 1438 994
rect 1382 956 1438 958
rect 1382 904 1384 956
rect 1384 904 1436 956
rect 1436 904 1438 956
rect 1382 902 1438 904
rect 1382 866 1438 868
rect 1382 814 1384 866
rect 1384 814 1436 866
rect 1436 814 1438 866
rect 1382 812 1438 814
rect 1682 1316 1738 1318
rect 1682 1264 1684 1316
rect 1684 1264 1736 1316
rect 1736 1264 1738 1316
rect 1682 1262 1738 1264
rect 1682 1226 1738 1228
rect 1682 1174 1684 1226
rect 1684 1174 1736 1226
rect 1736 1174 1738 1226
rect 1682 1172 1738 1174
rect 1682 1136 1738 1138
rect 1682 1084 1684 1136
rect 1684 1084 1736 1136
rect 1736 1084 1738 1136
rect 1682 1082 1738 1084
rect 1682 1046 1738 1048
rect 1682 994 1684 1046
rect 1684 994 1736 1046
rect 1736 994 1738 1046
rect 1682 992 1738 994
rect 1682 956 1738 958
rect 1682 904 1684 956
rect 1684 904 1736 956
rect 1736 904 1738 956
rect 1682 902 1738 904
rect 1682 866 1738 868
rect 1682 814 1684 866
rect 1684 814 1736 866
rect 1736 814 1738 866
rect 1682 812 1738 814
rect 1982 1316 2038 1318
rect 1982 1264 1984 1316
rect 1984 1264 2036 1316
rect 2036 1264 2038 1316
rect 1982 1262 2038 1264
rect 1982 1226 2038 1228
rect 1982 1174 1984 1226
rect 1984 1174 2036 1226
rect 2036 1174 2038 1226
rect 1982 1172 2038 1174
rect 1982 1136 2038 1138
rect 1982 1084 1984 1136
rect 1984 1084 2036 1136
rect 2036 1084 2038 1136
rect 1982 1082 2038 1084
rect 1982 1046 2038 1048
rect 1982 994 1984 1046
rect 1984 994 2036 1046
rect 2036 994 2038 1046
rect 1982 992 2038 994
rect 1982 956 2038 958
rect 1982 904 1984 956
rect 1984 904 2036 956
rect 2036 904 2038 956
rect 1982 902 2038 904
rect 1982 866 2038 868
rect 1982 814 1984 866
rect 1984 814 2036 866
rect 2036 814 2038 866
rect 1982 812 2038 814
rect 2282 1316 2338 1318
rect 2282 1264 2284 1316
rect 2284 1264 2336 1316
rect 2336 1264 2338 1316
rect 2282 1262 2338 1264
rect 2282 1226 2338 1228
rect 2282 1174 2284 1226
rect 2284 1174 2336 1226
rect 2336 1174 2338 1226
rect 2282 1172 2338 1174
rect 2282 1136 2338 1138
rect 2282 1084 2284 1136
rect 2284 1084 2336 1136
rect 2336 1084 2338 1136
rect 2282 1082 2338 1084
rect 2282 1046 2338 1048
rect 2282 994 2284 1046
rect 2284 994 2336 1046
rect 2336 994 2338 1046
rect 2282 992 2338 994
rect 2282 956 2338 958
rect 2282 904 2284 956
rect 2284 904 2336 956
rect 2336 904 2338 956
rect 2282 902 2338 904
rect 2282 866 2338 868
rect 2282 814 2284 866
rect 2284 814 2336 866
rect 2336 814 2338 866
rect 2282 812 2338 814
rect 2582 1316 2638 1318
rect 2582 1264 2584 1316
rect 2584 1264 2636 1316
rect 2636 1264 2638 1316
rect 2582 1262 2638 1264
rect 2582 1226 2638 1228
rect 2582 1174 2584 1226
rect 2584 1174 2636 1226
rect 2636 1174 2638 1226
rect 2582 1172 2638 1174
rect 2582 1136 2638 1138
rect 2582 1084 2584 1136
rect 2584 1084 2636 1136
rect 2636 1084 2638 1136
rect 2582 1082 2638 1084
rect 2582 1046 2638 1048
rect 2582 994 2584 1046
rect 2584 994 2636 1046
rect 2636 994 2638 1046
rect 2582 992 2638 994
rect 2582 956 2638 958
rect 2582 904 2584 956
rect 2584 904 2636 956
rect 2636 904 2638 956
rect 2582 902 2638 904
rect 2582 866 2638 868
rect 2582 814 2584 866
rect 2584 814 2636 866
rect 2636 814 2638 866
rect 2582 812 2638 814
rect 2882 1316 2938 1318
rect 2882 1264 2884 1316
rect 2884 1264 2936 1316
rect 2936 1264 2938 1316
rect 2882 1262 2938 1264
rect 2882 1226 2938 1228
rect 2882 1174 2884 1226
rect 2884 1174 2936 1226
rect 2936 1174 2938 1226
rect 2882 1172 2938 1174
rect 2882 1136 2938 1138
rect 2882 1084 2884 1136
rect 2884 1084 2936 1136
rect 2936 1084 2938 1136
rect 2882 1082 2938 1084
rect 2882 1046 2938 1048
rect 2882 994 2884 1046
rect 2884 994 2936 1046
rect 2936 994 2938 1046
rect 2882 992 2938 994
rect 2882 956 2938 958
rect 2882 904 2884 956
rect 2884 904 2936 956
rect 2936 904 2938 956
rect 2882 902 2938 904
rect 2882 866 2938 868
rect 2882 814 2884 866
rect 2884 814 2936 866
rect 2936 814 2938 866
rect 2882 812 2938 814
rect 3482 1316 3538 1318
rect 3482 1264 3484 1316
rect 3484 1264 3536 1316
rect 3536 1264 3538 1316
rect 3482 1262 3538 1264
rect 3482 1226 3538 1228
rect 3482 1174 3484 1226
rect 3484 1174 3536 1226
rect 3536 1174 3538 1226
rect 3482 1172 3538 1174
rect 3482 1136 3538 1138
rect 3482 1084 3484 1136
rect 3484 1084 3536 1136
rect 3536 1084 3538 1136
rect 3482 1082 3538 1084
rect 3482 1046 3538 1048
rect 3482 994 3484 1046
rect 3484 994 3536 1046
rect 3536 994 3538 1046
rect 3482 992 3538 994
rect 3482 956 3538 958
rect 3482 904 3484 956
rect 3484 904 3536 956
rect 3536 904 3538 956
rect 3482 902 3538 904
rect 3482 866 3538 868
rect 3482 814 3484 866
rect 3484 814 3536 866
rect 3536 814 3538 866
rect 3482 812 3538 814
rect 3782 1316 3838 1318
rect 3782 1264 3784 1316
rect 3784 1264 3836 1316
rect 3836 1264 3838 1316
rect 3782 1262 3838 1264
rect 3782 1226 3838 1228
rect 3782 1174 3784 1226
rect 3784 1174 3836 1226
rect 3836 1174 3838 1226
rect 3782 1172 3838 1174
rect 3782 1136 3838 1138
rect 3782 1084 3784 1136
rect 3784 1084 3836 1136
rect 3836 1084 3838 1136
rect 3782 1082 3838 1084
rect 3782 1046 3838 1048
rect 3782 994 3784 1046
rect 3784 994 3836 1046
rect 3836 994 3838 1046
rect 3782 992 3838 994
rect 3782 956 3838 958
rect 3782 904 3784 956
rect 3784 904 3836 956
rect 3836 904 3838 956
rect 3782 902 3838 904
rect 3782 866 3838 868
rect 3782 814 3784 866
rect 3784 814 3836 866
rect 3836 814 3838 866
rect 3782 812 3838 814
rect 4082 1316 4138 1318
rect 4082 1264 4084 1316
rect 4084 1264 4136 1316
rect 4136 1264 4138 1316
rect 4082 1262 4138 1264
rect 4082 1226 4138 1228
rect 4082 1174 4084 1226
rect 4084 1174 4136 1226
rect 4136 1174 4138 1226
rect 4082 1172 4138 1174
rect 4082 1136 4138 1138
rect 4082 1084 4084 1136
rect 4084 1084 4136 1136
rect 4136 1084 4138 1136
rect 4082 1082 4138 1084
rect 4082 1046 4138 1048
rect 4082 994 4084 1046
rect 4084 994 4136 1046
rect 4136 994 4138 1046
rect 4082 992 4138 994
rect 4082 956 4138 958
rect 4082 904 4084 956
rect 4084 904 4136 956
rect 4136 904 4138 956
rect 4082 902 4138 904
rect 4082 866 4138 868
rect 4082 814 4084 866
rect 4084 814 4136 866
rect 4136 814 4138 866
rect 4082 812 4138 814
rect 4382 1316 4438 1318
rect 4382 1264 4384 1316
rect 4384 1264 4436 1316
rect 4436 1264 4438 1316
rect 4382 1262 4438 1264
rect 4382 1226 4438 1228
rect 4382 1174 4384 1226
rect 4384 1174 4436 1226
rect 4436 1174 4438 1226
rect 4382 1172 4438 1174
rect 4382 1136 4438 1138
rect 4382 1084 4384 1136
rect 4384 1084 4436 1136
rect 4436 1084 4438 1136
rect 4382 1082 4438 1084
rect 4382 1046 4438 1048
rect 4382 994 4384 1046
rect 4384 994 4436 1046
rect 4436 994 4438 1046
rect 4382 992 4438 994
rect 4382 956 4438 958
rect 4382 904 4384 956
rect 4384 904 4436 956
rect 4436 904 4438 956
rect 4382 902 4438 904
rect 4382 866 4438 868
rect 4382 814 4384 866
rect 4384 814 4436 866
rect 4436 814 4438 866
rect 4382 812 4438 814
rect 4682 1316 4738 1318
rect 4682 1264 4684 1316
rect 4684 1264 4736 1316
rect 4736 1264 4738 1316
rect 4682 1262 4738 1264
rect 4682 1226 4738 1228
rect 4682 1174 4684 1226
rect 4684 1174 4736 1226
rect 4736 1174 4738 1226
rect 4682 1172 4738 1174
rect 4682 1136 4738 1138
rect 4682 1084 4684 1136
rect 4684 1084 4736 1136
rect 4736 1084 4738 1136
rect 4682 1082 4738 1084
rect 4682 1046 4738 1048
rect 4682 994 4684 1046
rect 4684 994 4736 1046
rect 4736 994 4738 1046
rect 4682 992 4738 994
rect 4682 956 4738 958
rect 4682 904 4684 956
rect 4684 904 4736 956
rect 4736 904 4738 956
rect 4682 902 4738 904
rect 4682 866 4738 868
rect 4682 814 4684 866
rect 4684 814 4736 866
rect 4736 814 4738 866
rect 4682 812 4738 814
rect 4982 1316 5038 1318
rect 4982 1264 4984 1316
rect 4984 1264 5036 1316
rect 5036 1264 5038 1316
rect 4982 1262 5038 1264
rect 4982 1226 5038 1228
rect 4982 1174 4984 1226
rect 4984 1174 5036 1226
rect 5036 1174 5038 1226
rect 4982 1172 5038 1174
rect 4982 1136 5038 1138
rect 4982 1084 4984 1136
rect 4984 1084 5036 1136
rect 5036 1084 5038 1136
rect 4982 1082 5038 1084
rect 4982 1046 5038 1048
rect 4982 994 4984 1046
rect 4984 994 5036 1046
rect 5036 994 5038 1046
rect 4982 992 5038 994
rect 4982 956 5038 958
rect 4982 904 4984 956
rect 4984 904 5036 956
rect 5036 904 5038 956
rect 4982 902 5038 904
rect 4982 866 5038 868
rect 4982 814 4984 866
rect 4984 814 5036 866
rect 5036 814 5038 866
rect 4982 812 5038 814
rect 5282 1316 5338 1318
rect 5282 1264 5284 1316
rect 5284 1264 5336 1316
rect 5336 1264 5338 1316
rect 5282 1262 5338 1264
rect 5282 1226 5338 1228
rect 5282 1174 5284 1226
rect 5284 1174 5336 1226
rect 5336 1174 5338 1226
rect 5282 1172 5338 1174
rect 5282 1136 5338 1138
rect 5282 1084 5284 1136
rect 5284 1084 5336 1136
rect 5336 1084 5338 1136
rect 5282 1082 5338 1084
rect 5282 1046 5338 1048
rect 5282 994 5284 1046
rect 5284 994 5336 1046
rect 5336 994 5338 1046
rect 5282 992 5338 994
rect 5282 956 5338 958
rect 5282 904 5284 956
rect 5284 904 5336 956
rect 5336 904 5338 956
rect 5282 902 5338 904
rect 5282 866 5338 868
rect 5282 814 5284 866
rect 5284 814 5336 866
rect 5336 814 5338 866
rect 5282 812 5338 814
rect 5582 1316 5638 1318
rect 5582 1264 5584 1316
rect 5584 1264 5636 1316
rect 5636 1264 5638 1316
rect 5582 1262 5638 1264
rect 5582 1226 5638 1228
rect 5582 1174 5584 1226
rect 5584 1174 5636 1226
rect 5636 1174 5638 1226
rect 5582 1172 5638 1174
rect 5582 1136 5638 1138
rect 5582 1084 5584 1136
rect 5584 1084 5636 1136
rect 5636 1084 5638 1136
rect 5582 1082 5638 1084
rect 5582 1046 5638 1048
rect 5582 994 5584 1046
rect 5584 994 5636 1046
rect 5636 994 5638 1046
rect 5582 992 5638 994
rect 5582 956 5638 958
rect 5582 904 5584 956
rect 5584 904 5636 956
rect 5636 904 5638 956
rect 5582 902 5638 904
rect 5582 866 5638 868
rect 5582 814 5584 866
rect 5584 814 5636 866
rect 5636 814 5638 866
rect 5582 812 5638 814
rect 5882 1316 5938 1318
rect 5882 1264 5884 1316
rect 5884 1264 5936 1316
rect 5936 1264 5938 1316
rect 5882 1262 5938 1264
rect 5882 1226 5938 1228
rect 5882 1174 5884 1226
rect 5884 1174 5936 1226
rect 5936 1174 5938 1226
rect 5882 1172 5938 1174
rect 5882 1136 5938 1138
rect 5882 1084 5884 1136
rect 5884 1084 5936 1136
rect 5936 1084 5938 1136
rect 5882 1082 5938 1084
rect 5882 1046 5938 1048
rect 5882 994 5884 1046
rect 5884 994 5936 1046
rect 5936 994 5938 1046
rect 5882 992 5938 994
rect 5882 956 5938 958
rect 5882 904 5884 956
rect 5884 904 5936 956
rect 5936 904 5938 956
rect 5882 902 5938 904
rect 5882 866 5938 868
rect 5882 814 5884 866
rect 5884 814 5936 866
rect 5936 814 5938 866
rect 5882 812 5938 814
rect 6182 1316 6238 1318
rect 6182 1264 6184 1316
rect 6184 1264 6236 1316
rect 6236 1264 6238 1316
rect 6182 1262 6238 1264
rect 6182 1226 6238 1228
rect 6182 1174 6184 1226
rect 6184 1174 6236 1226
rect 6236 1174 6238 1226
rect 6182 1172 6238 1174
rect 6182 1136 6238 1138
rect 6182 1084 6184 1136
rect 6184 1084 6236 1136
rect 6236 1084 6238 1136
rect 6182 1082 6238 1084
rect 6182 1046 6238 1048
rect 6182 994 6184 1046
rect 6184 994 6236 1046
rect 6236 994 6238 1046
rect 6182 992 6238 994
rect 6182 956 6238 958
rect 6182 904 6184 956
rect 6184 904 6236 956
rect 6236 904 6238 956
rect 6182 902 6238 904
rect 6182 866 6238 868
rect 6182 814 6184 866
rect 6184 814 6236 866
rect 6236 814 6238 866
rect 6182 812 6238 814
rect -58 142 -2 198
rect -198 52 -142 108
rect -58 52 -2 108
rect 6582 142 6638 198
rect 6582 52 6638 108
rect 6722 52 6778 108
rect -198 -38 -142 18
rect 6722 -38 6778 18
rect -58 -278 -2 -222
rect -198 -368 -142 -312
rect -58 -368 -2 -312
rect 6582 -278 6638 -222
rect 6582 -368 6638 -312
rect 6722 -368 6778 -312
rect -198 -458 -142 -402
rect 6722 -458 6778 -402
<< metal3 >>
rect 6467 5268 6577 5290
rect 6467 5212 6494 5268
rect 6550 5212 6577 5268
rect 6467 5190 6577 5212
rect 6707 5268 6817 5290
rect 6707 5212 6734 5268
rect 6790 5212 6817 5268
rect 6707 5190 6817 5212
rect 470 5042 570 5060
rect 470 4978 488 5042
rect 552 4978 570 5042
rect 470 4960 570 4978
rect 770 5042 870 5060
rect 770 4978 788 5042
rect 852 4978 870 5042
rect 770 4960 870 4978
rect 1070 5042 1170 5060
rect 1070 4978 1088 5042
rect 1152 4978 1170 5042
rect 1070 4960 1170 4978
rect 1370 5042 1470 5060
rect 1370 4978 1388 5042
rect 1452 4978 1470 5042
rect 1370 4960 1470 4978
rect 1670 5042 1770 5060
rect 1670 4978 1688 5042
rect 1752 4978 1770 5042
rect 1670 4960 1770 4978
rect 1970 5042 2070 5060
rect 1970 4978 1988 5042
rect 2052 4978 2070 5042
rect 1970 4960 2070 4978
rect 2270 5042 2370 5060
rect 2270 4978 2288 5042
rect 2352 4978 2370 5042
rect 2270 4960 2370 4978
rect 2570 5042 2670 5060
rect 2570 4978 2588 5042
rect 2652 4978 2670 5042
rect 2570 4960 2670 4978
rect 2870 5042 2970 5060
rect 2870 4978 2888 5042
rect 2952 4978 2970 5042
rect 2870 4960 2970 4978
rect 3170 5042 3270 5060
rect 3170 4978 3188 5042
rect 3252 4978 3270 5042
rect 3170 4960 3270 4978
rect 3470 5042 3570 5060
rect 3470 4978 3488 5042
rect 3552 4978 3570 5042
rect 3470 4960 3570 4978
rect 3770 5042 3870 5060
rect 3770 4978 3788 5042
rect 3852 4978 3870 5042
rect 3770 4960 3870 4978
rect 4070 5042 4170 5060
rect 4070 4978 4088 5042
rect 4152 4978 4170 5042
rect 4070 4960 4170 4978
rect 4370 5042 4470 5060
rect 4370 4978 4388 5042
rect 4452 4978 4470 5042
rect 4370 4960 4470 4978
rect 4670 5042 4770 5060
rect 4670 4978 4688 5042
rect 4752 4978 4770 5042
rect 4670 4960 4770 4978
rect 4970 5042 5070 5060
rect 4970 4978 4988 5042
rect 5052 4978 5070 5042
rect 4970 4960 5070 4978
rect 5270 5042 5370 5060
rect 5270 4978 5288 5042
rect 5352 4978 5370 5042
rect 5270 4960 5370 4978
rect 5570 5042 5670 5060
rect 5570 4978 5588 5042
rect 5652 4978 5670 5042
rect 5570 4960 5670 4978
rect 5870 5042 5970 5060
rect 5870 4978 5888 5042
rect 5952 4978 5970 5042
rect 5870 4960 5970 4978
rect 6170 5042 6270 5060
rect 6170 4978 6188 5042
rect 6252 4978 6270 5042
rect 6170 4960 6270 4978
rect 490 3650 550 4960
rect 790 3650 850 4960
rect 1090 3650 1150 4960
rect 1390 3650 1450 4960
rect 1690 3650 1750 4960
rect 1990 3650 2050 4960
rect 2290 3650 2350 4960
rect 2590 3650 2650 4960
rect 2890 3650 2950 4960
rect 3190 3650 3250 4960
rect 470 3628 550 3650
rect 470 3572 482 3628
rect 538 3572 550 3628
rect 470 3538 550 3572
rect 470 3482 482 3538
rect 538 3482 550 3538
rect 470 3448 550 3482
rect 470 3392 482 3448
rect 538 3392 550 3448
rect 470 3358 550 3392
rect 470 3302 482 3358
rect 538 3302 550 3358
rect 470 3268 550 3302
rect 470 3212 482 3268
rect 538 3212 550 3268
rect 470 3178 550 3212
rect 470 3122 482 3178
rect 538 3122 550 3178
rect 470 3110 550 3122
rect 770 3628 850 3650
rect 770 3572 782 3628
rect 838 3572 850 3628
rect 770 3538 850 3572
rect 770 3482 782 3538
rect 838 3482 850 3538
rect 770 3448 850 3482
rect 770 3392 782 3448
rect 838 3392 850 3448
rect 770 3358 850 3392
rect 770 3302 782 3358
rect 838 3302 850 3358
rect 770 3268 850 3302
rect 770 3212 782 3268
rect 838 3212 850 3268
rect 770 3178 850 3212
rect 770 3122 782 3178
rect 838 3122 850 3178
rect 770 3110 850 3122
rect 1070 3628 1150 3650
rect 1070 3572 1082 3628
rect 1138 3572 1150 3628
rect 1070 3538 1150 3572
rect 1070 3482 1082 3538
rect 1138 3482 1150 3538
rect 1070 3448 1150 3482
rect 1070 3392 1082 3448
rect 1138 3392 1150 3448
rect 1070 3358 1150 3392
rect 1070 3302 1082 3358
rect 1138 3302 1150 3358
rect 1070 3268 1150 3302
rect 1070 3212 1082 3268
rect 1138 3212 1150 3268
rect 1070 3178 1150 3212
rect 1070 3122 1082 3178
rect 1138 3122 1150 3178
rect 1070 3110 1150 3122
rect 1370 3628 1450 3650
rect 1370 3572 1382 3628
rect 1438 3572 1450 3628
rect 1370 3538 1450 3572
rect 1370 3482 1382 3538
rect 1438 3482 1450 3538
rect 1370 3448 1450 3482
rect 1370 3392 1382 3448
rect 1438 3392 1450 3448
rect 1370 3358 1450 3392
rect 1370 3302 1382 3358
rect 1438 3302 1450 3358
rect 1370 3268 1450 3302
rect 1370 3212 1382 3268
rect 1438 3212 1450 3268
rect 1370 3178 1450 3212
rect 1370 3122 1382 3178
rect 1438 3122 1450 3178
rect 1370 3110 1450 3122
rect 1670 3628 1750 3650
rect 1670 3572 1682 3628
rect 1738 3572 1750 3628
rect 1670 3538 1750 3572
rect 1670 3482 1682 3538
rect 1738 3482 1750 3538
rect 1670 3448 1750 3482
rect 1670 3392 1682 3448
rect 1738 3392 1750 3448
rect 1670 3358 1750 3392
rect 1670 3302 1682 3358
rect 1738 3302 1750 3358
rect 1670 3268 1750 3302
rect 1670 3212 1682 3268
rect 1738 3212 1750 3268
rect 1670 3178 1750 3212
rect 1670 3122 1682 3178
rect 1738 3122 1750 3178
rect 1670 3110 1750 3122
rect 1970 3628 2050 3650
rect 1970 3572 1982 3628
rect 2038 3572 2050 3628
rect 1970 3538 2050 3572
rect 1970 3482 1982 3538
rect 2038 3482 2050 3538
rect 1970 3448 2050 3482
rect 1970 3392 1982 3448
rect 2038 3392 2050 3448
rect 1970 3358 2050 3392
rect 1970 3302 1982 3358
rect 2038 3302 2050 3358
rect 1970 3268 2050 3302
rect 1970 3212 1982 3268
rect 2038 3212 2050 3268
rect 1970 3178 2050 3212
rect 1970 3122 1982 3178
rect 2038 3122 2050 3178
rect 1970 3110 2050 3122
rect 2270 3628 2350 3650
rect 2270 3572 2282 3628
rect 2338 3572 2350 3628
rect 2270 3538 2350 3572
rect 2270 3482 2282 3538
rect 2338 3482 2350 3538
rect 2270 3448 2350 3482
rect 2270 3392 2282 3448
rect 2338 3392 2350 3448
rect 2270 3358 2350 3392
rect 2270 3302 2282 3358
rect 2338 3302 2350 3358
rect 2270 3268 2350 3302
rect 2270 3212 2282 3268
rect 2338 3212 2350 3268
rect 2270 3178 2350 3212
rect 2270 3122 2282 3178
rect 2338 3122 2350 3178
rect 2270 3110 2350 3122
rect 2570 3628 2650 3650
rect 2570 3572 2582 3628
rect 2638 3572 2650 3628
rect 2570 3538 2650 3572
rect 2570 3482 2582 3538
rect 2638 3482 2650 3538
rect 2570 3448 2650 3482
rect 2570 3392 2582 3448
rect 2638 3392 2650 3448
rect 2570 3358 2650 3392
rect 2570 3302 2582 3358
rect 2638 3302 2650 3358
rect 2570 3268 2650 3302
rect 2570 3212 2582 3268
rect 2638 3212 2650 3268
rect 2570 3178 2650 3212
rect 2570 3122 2582 3178
rect 2638 3122 2650 3178
rect 2570 3110 2650 3122
rect 2870 3628 2950 3650
rect 2870 3572 2882 3628
rect 2938 3572 2950 3628
rect 2870 3538 2950 3572
rect 2870 3482 2882 3538
rect 2938 3482 2950 3538
rect 2870 3448 2950 3482
rect 2870 3392 2882 3448
rect 2938 3392 2950 3448
rect 2870 3358 2950 3392
rect 2870 3302 2882 3358
rect 2938 3302 2950 3358
rect 2870 3268 2950 3302
rect 2870 3212 2882 3268
rect 2938 3212 2950 3268
rect 2870 3178 2950 3212
rect 2870 3122 2882 3178
rect 2938 3122 2950 3178
rect 2870 3110 2950 3122
rect 3170 3628 3250 3650
rect 3170 3572 3182 3628
rect 3238 3572 3250 3628
rect 3170 3538 3250 3572
rect 3170 3482 3182 3538
rect 3238 3482 3250 3538
rect 3170 3448 3250 3482
rect 3170 3392 3182 3448
rect 3238 3392 3250 3448
rect 3170 3358 3250 3392
rect 3170 3302 3182 3358
rect 3238 3302 3250 3358
rect 3170 3268 3250 3302
rect 3170 3212 3182 3268
rect 3238 3212 3250 3268
rect 3170 3178 3250 3212
rect 3170 3122 3182 3178
rect 3238 3122 3250 3178
rect 3170 3110 3250 3122
rect -70 2518 10 2530
rect -70 2462 -58 2518
rect -2 2462 10 2518
rect -210 2428 -130 2440
rect -210 2372 -198 2428
rect -142 2372 -130 2428
rect -210 2338 -130 2372
rect -210 2282 -198 2338
rect -142 2282 -130 2338
rect -210 108 -130 2282
rect -210 52 -198 108
rect -142 52 -130 108
rect -210 18 -130 52
rect -210 -38 -198 18
rect -142 -38 -130 18
rect -210 -312 -130 -38
rect -210 -368 -198 -312
rect -142 -368 -130 -312
rect -210 -402 -130 -368
rect -70 2428 10 2462
rect -70 2372 -58 2428
rect -2 2372 10 2428
rect -70 198 10 2372
rect 490 1340 550 3110
rect 790 1340 850 3110
rect 1090 1340 1150 3110
rect 1390 1340 1450 3110
rect 1690 1340 1750 3110
rect 1990 1340 2050 3110
rect 2290 1340 2350 3110
rect 2590 1340 2650 3110
rect 2890 1340 2950 3110
rect 3190 2710 3250 3110
rect 3490 1340 3550 4960
rect 3790 3650 3850 4960
rect 4090 3650 4150 4960
rect 4390 3650 4450 4960
rect 4690 3650 4750 4960
rect 4990 3650 5050 4960
rect 5290 3650 5350 4960
rect 5590 3650 5650 4960
rect 5890 3650 5950 4960
rect 6190 3650 6250 4960
rect 3770 3628 3850 3650
rect 3770 3572 3782 3628
rect 3838 3572 3850 3628
rect 3770 3538 3850 3572
rect 3770 3482 3782 3538
rect 3838 3482 3850 3538
rect 3770 3448 3850 3482
rect 3770 3392 3782 3448
rect 3838 3392 3850 3448
rect 3770 3358 3850 3392
rect 3770 3302 3782 3358
rect 3838 3302 3850 3358
rect 3770 3268 3850 3302
rect 3770 3212 3782 3268
rect 3838 3212 3850 3268
rect 3770 3178 3850 3212
rect 3770 3122 3782 3178
rect 3838 3122 3850 3178
rect 3770 3110 3850 3122
rect 4070 3628 4150 3650
rect 4070 3572 4082 3628
rect 4138 3572 4150 3628
rect 4070 3538 4150 3572
rect 4070 3482 4082 3538
rect 4138 3482 4150 3538
rect 4070 3448 4150 3482
rect 4070 3392 4082 3448
rect 4138 3392 4150 3448
rect 4070 3358 4150 3392
rect 4070 3302 4082 3358
rect 4138 3302 4150 3358
rect 4070 3268 4150 3302
rect 4070 3212 4082 3268
rect 4138 3212 4150 3268
rect 4070 3178 4150 3212
rect 4070 3122 4082 3178
rect 4138 3122 4150 3178
rect 4070 3110 4150 3122
rect 4370 3628 4450 3650
rect 4370 3572 4382 3628
rect 4438 3572 4450 3628
rect 4370 3538 4450 3572
rect 4370 3482 4382 3538
rect 4438 3482 4450 3538
rect 4370 3448 4450 3482
rect 4370 3392 4382 3448
rect 4438 3392 4450 3448
rect 4370 3358 4450 3392
rect 4370 3302 4382 3358
rect 4438 3302 4450 3358
rect 4370 3268 4450 3302
rect 4370 3212 4382 3268
rect 4438 3212 4450 3268
rect 4370 3178 4450 3212
rect 4370 3122 4382 3178
rect 4438 3122 4450 3178
rect 4370 3110 4450 3122
rect 4670 3628 4750 3650
rect 4670 3572 4682 3628
rect 4738 3572 4750 3628
rect 4670 3538 4750 3572
rect 4670 3482 4682 3538
rect 4738 3482 4750 3538
rect 4670 3448 4750 3482
rect 4670 3392 4682 3448
rect 4738 3392 4750 3448
rect 4670 3358 4750 3392
rect 4670 3302 4682 3358
rect 4738 3302 4750 3358
rect 4670 3268 4750 3302
rect 4670 3212 4682 3268
rect 4738 3212 4750 3268
rect 4670 3178 4750 3212
rect 4670 3122 4682 3178
rect 4738 3122 4750 3178
rect 4670 3110 4750 3122
rect 4970 3628 5050 3650
rect 4970 3572 4982 3628
rect 5038 3572 5050 3628
rect 4970 3538 5050 3572
rect 4970 3482 4982 3538
rect 5038 3482 5050 3538
rect 4970 3448 5050 3482
rect 4970 3392 4982 3448
rect 5038 3392 5050 3448
rect 4970 3358 5050 3392
rect 4970 3302 4982 3358
rect 5038 3302 5050 3358
rect 4970 3268 5050 3302
rect 4970 3212 4982 3268
rect 5038 3212 5050 3268
rect 4970 3178 5050 3212
rect 4970 3122 4982 3178
rect 5038 3122 5050 3178
rect 4970 3110 5050 3122
rect 5270 3628 5350 3650
rect 5270 3572 5282 3628
rect 5338 3572 5350 3628
rect 5270 3538 5350 3572
rect 5270 3482 5282 3538
rect 5338 3482 5350 3538
rect 5270 3448 5350 3482
rect 5270 3392 5282 3448
rect 5338 3392 5350 3448
rect 5270 3358 5350 3392
rect 5270 3302 5282 3358
rect 5338 3302 5350 3358
rect 5270 3268 5350 3302
rect 5270 3212 5282 3268
rect 5338 3212 5350 3268
rect 5270 3178 5350 3212
rect 5270 3122 5282 3178
rect 5338 3122 5350 3178
rect 5270 3110 5350 3122
rect 5570 3628 5650 3650
rect 5570 3572 5582 3628
rect 5638 3572 5650 3628
rect 5570 3538 5650 3572
rect 5570 3482 5582 3538
rect 5638 3482 5650 3538
rect 5570 3448 5650 3482
rect 5570 3392 5582 3448
rect 5638 3392 5650 3448
rect 5570 3358 5650 3392
rect 5570 3302 5582 3358
rect 5638 3302 5650 3358
rect 5570 3268 5650 3302
rect 5570 3212 5582 3268
rect 5638 3212 5650 3268
rect 5570 3178 5650 3212
rect 5570 3122 5582 3178
rect 5638 3122 5650 3178
rect 5570 3110 5650 3122
rect 5870 3628 5950 3650
rect 5870 3572 5882 3628
rect 5938 3572 5950 3628
rect 5870 3538 5950 3572
rect 5870 3482 5882 3538
rect 5938 3482 5950 3538
rect 5870 3448 5950 3482
rect 5870 3392 5882 3448
rect 5938 3392 5950 3448
rect 5870 3358 5950 3392
rect 5870 3302 5882 3358
rect 5938 3302 5950 3358
rect 5870 3268 5950 3302
rect 5870 3212 5882 3268
rect 5938 3212 5950 3268
rect 5870 3178 5950 3212
rect 5870 3122 5882 3178
rect 5938 3122 5950 3178
rect 5870 3110 5950 3122
rect 6170 3628 6250 3650
rect 6170 3572 6182 3628
rect 6238 3572 6250 3628
rect 6170 3538 6250 3572
rect 6170 3482 6182 3538
rect 6238 3482 6250 3538
rect 6170 3448 6250 3482
rect 6170 3392 6182 3448
rect 6238 3392 6250 3448
rect 6170 3358 6250 3392
rect 6170 3302 6182 3358
rect 6238 3302 6250 3358
rect 6170 3268 6250 3302
rect 6170 3212 6182 3268
rect 6238 3212 6250 3268
rect 6170 3178 6250 3212
rect 6170 3122 6182 3178
rect 6238 3122 6250 3178
rect 6170 3110 6250 3122
rect 3790 1340 3850 3110
rect 4090 1340 4150 3110
rect 4390 1340 4450 3110
rect 4690 1340 4750 3110
rect 4990 1340 5050 3110
rect 5290 1340 5350 3110
rect 5590 1340 5650 3110
rect 5890 1340 5950 3110
rect 6190 1340 6250 3110
rect 470 1318 550 1340
rect 470 1262 482 1318
rect 538 1262 550 1318
rect 470 1228 550 1262
rect 470 1172 482 1228
rect 538 1172 550 1228
rect 470 1138 550 1172
rect 470 1082 482 1138
rect 538 1082 550 1138
rect 470 1048 550 1082
rect 470 992 482 1048
rect 538 992 550 1048
rect 470 958 550 992
rect 470 902 482 958
rect 538 902 550 958
rect 470 868 550 902
rect 470 812 482 868
rect 538 812 550 868
rect 470 800 550 812
rect 770 1318 850 1340
rect 770 1262 782 1318
rect 838 1262 850 1318
rect 770 1228 850 1262
rect 770 1172 782 1228
rect 838 1172 850 1228
rect 770 1138 850 1172
rect 770 1082 782 1138
rect 838 1082 850 1138
rect 770 1048 850 1082
rect 770 992 782 1048
rect 838 992 850 1048
rect 770 958 850 992
rect 770 902 782 958
rect 838 902 850 958
rect 770 868 850 902
rect 770 812 782 868
rect 838 812 850 868
rect 770 800 850 812
rect 1070 1318 1150 1340
rect 1070 1262 1082 1318
rect 1138 1262 1150 1318
rect 1070 1228 1150 1262
rect 1070 1172 1082 1228
rect 1138 1172 1150 1228
rect 1070 1138 1150 1172
rect 1070 1082 1082 1138
rect 1138 1082 1150 1138
rect 1070 1048 1150 1082
rect 1070 992 1082 1048
rect 1138 992 1150 1048
rect 1070 958 1150 992
rect 1070 902 1082 958
rect 1138 902 1150 958
rect 1070 868 1150 902
rect 1070 812 1082 868
rect 1138 812 1150 868
rect 1070 800 1150 812
rect 1370 1318 1450 1340
rect 1370 1262 1382 1318
rect 1438 1262 1450 1318
rect 1370 1228 1450 1262
rect 1370 1172 1382 1228
rect 1438 1172 1450 1228
rect 1370 1138 1450 1172
rect 1370 1082 1382 1138
rect 1438 1082 1450 1138
rect 1370 1048 1450 1082
rect 1370 992 1382 1048
rect 1438 992 1450 1048
rect 1370 958 1450 992
rect 1370 902 1382 958
rect 1438 902 1450 958
rect 1370 868 1450 902
rect 1370 812 1382 868
rect 1438 812 1450 868
rect 1370 800 1450 812
rect 1670 1318 1750 1340
rect 1670 1262 1682 1318
rect 1738 1262 1750 1318
rect 1670 1228 1750 1262
rect 1670 1172 1682 1228
rect 1738 1172 1750 1228
rect 1670 1138 1750 1172
rect 1670 1082 1682 1138
rect 1738 1082 1750 1138
rect 1670 1048 1750 1082
rect 1670 992 1682 1048
rect 1738 992 1750 1048
rect 1670 958 1750 992
rect 1670 902 1682 958
rect 1738 902 1750 958
rect 1670 868 1750 902
rect 1670 812 1682 868
rect 1738 812 1750 868
rect 1670 800 1750 812
rect 1970 1318 2050 1340
rect 1970 1262 1982 1318
rect 2038 1262 2050 1318
rect 1970 1228 2050 1262
rect 1970 1172 1982 1228
rect 2038 1172 2050 1228
rect 1970 1138 2050 1172
rect 1970 1082 1982 1138
rect 2038 1082 2050 1138
rect 1970 1048 2050 1082
rect 1970 992 1982 1048
rect 2038 992 2050 1048
rect 1970 958 2050 992
rect 1970 902 1982 958
rect 2038 902 2050 958
rect 1970 868 2050 902
rect 1970 812 1982 868
rect 2038 812 2050 868
rect 1970 800 2050 812
rect 2270 1318 2350 1340
rect 2270 1262 2282 1318
rect 2338 1262 2350 1318
rect 2270 1228 2350 1262
rect 2270 1172 2282 1228
rect 2338 1172 2350 1228
rect 2270 1138 2350 1172
rect 2270 1082 2282 1138
rect 2338 1082 2350 1138
rect 2270 1048 2350 1082
rect 2270 992 2282 1048
rect 2338 992 2350 1048
rect 2270 958 2350 992
rect 2270 902 2282 958
rect 2338 902 2350 958
rect 2270 868 2350 902
rect 2270 812 2282 868
rect 2338 812 2350 868
rect 2270 800 2350 812
rect 2570 1318 2650 1340
rect 2570 1262 2582 1318
rect 2638 1262 2650 1318
rect 2570 1228 2650 1262
rect 2570 1172 2582 1228
rect 2638 1172 2650 1228
rect 2570 1138 2650 1172
rect 2570 1082 2582 1138
rect 2638 1082 2650 1138
rect 2570 1048 2650 1082
rect 2570 992 2582 1048
rect 2638 992 2650 1048
rect 2570 958 2650 992
rect 2570 902 2582 958
rect 2638 902 2650 958
rect 2570 868 2650 902
rect 2570 812 2582 868
rect 2638 812 2650 868
rect 2570 800 2650 812
rect 2870 1318 2950 1340
rect 2870 1262 2882 1318
rect 2938 1262 2950 1318
rect 2870 1228 2950 1262
rect 2870 1172 2882 1228
rect 2938 1172 2950 1228
rect 2870 1138 2950 1172
rect 2870 1082 2882 1138
rect 2938 1082 2950 1138
rect 2870 1048 2950 1082
rect 2870 992 2882 1048
rect 2938 992 2950 1048
rect 2870 958 2950 992
rect 2870 902 2882 958
rect 2938 902 2950 958
rect 2870 868 2950 902
rect 2870 812 2882 868
rect 2938 812 2950 868
rect 2870 800 2950 812
rect 3470 1318 3550 1340
rect 3470 1262 3482 1318
rect 3538 1262 3550 1318
rect 3470 1228 3550 1262
rect 3470 1172 3482 1228
rect 3538 1172 3550 1228
rect 3470 1138 3550 1172
rect 3470 1082 3482 1138
rect 3538 1082 3550 1138
rect 3470 1048 3550 1082
rect 3470 992 3482 1048
rect 3538 992 3550 1048
rect 3470 958 3550 992
rect 3470 902 3482 958
rect 3538 902 3550 958
rect 3470 868 3550 902
rect 3470 812 3482 868
rect 3538 812 3550 868
rect 3470 800 3550 812
rect 3770 1318 3850 1340
rect 3770 1262 3782 1318
rect 3838 1262 3850 1318
rect 3770 1228 3850 1262
rect 3770 1172 3782 1228
rect 3838 1172 3850 1228
rect 3770 1138 3850 1172
rect 3770 1082 3782 1138
rect 3838 1082 3850 1138
rect 3770 1048 3850 1082
rect 3770 992 3782 1048
rect 3838 992 3850 1048
rect 3770 958 3850 992
rect 3770 902 3782 958
rect 3838 902 3850 958
rect 3770 868 3850 902
rect 3770 812 3782 868
rect 3838 812 3850 868
rect 3770 800 3850 812
rect 4070 1318 4150 1340
rect 4070 1262 4082 1318
rect 4138 1262 4150 1318
rect 4070 1228 4150 1262
rect 4070 1172 4082 1228
rect 4138 1172 4150 1228
rect 4070 1138 4150 1172
rect 4070 1082 4082 1138
rect 4138 1082 4150 1138
rect 4070 1048 4150 1082
rect 4070 992 4082 1048
rect 4138 992 4150 1048
rect 4070 958 4150 992
rect 4070 902 4082 958
rect 4138 902 4150 958
rect 4070 868 4150 902
rect 4070 812 4082 868
rect 4138 812 4150 868
rect 4070 800 4150 812
rect 4370 1318 4450 1340
rect 4370 1262 4382 1318
rect 4438 1262 4450 1318
rect 4370 1228 4450 1262
rect 4370 1172 4382 1228
rect 4438 1172 4450 1228
rect 4370 1138 4450 1172
rect 4370 1082 4382 1138
rect 4438 1082 4450 1138
rect 4370 1048 4450 1082
rect 4370 992 4382 1048
rect 4438 992 4450 1048
rect 4370 958 4450 992
rect 4370 902 4382 958
rect 4438 902 4450 958
rect 4370 868 4450 902
rect 4370 812 4382 868
rect 4438 812 4450 868
rect 4370 800 4450 812
rect 4670 1318 4750 1340
rect 4670 1262 4682 1318
rect 4738 1262 4750 1318
rect 4670 1228 4750 1262
rect 4670 1172 4682 1228
rect 4738 1172 4750 1228
rect 4670 1138 4750 1172
rect 4670 1082 4682 1138
rect 4738 1082 4750 1138
rect 4670 1048 4750 1082
rect 4670 992 4682 1048
rect 4738 992 4750 1048
rect 4670 958 4750 992
rect 4670 902 4682 958
rect 4738 902 4750 958
rect 4670 868 4750 902
rect 4670 812 4682 868
rect 4738 812 4750 868
rect 4670 800 4750 812
rect 4970 1318 5050 1340
rect 4970 1262 4982 1318
rect 5038 1262 5050 1318
rect 4970 1228 5050 1262
rect 4970 1172 4982 1228
rect 5038 1172 5050 1228
rect 4970 1138 5050 1172
rect 4970 1082 4982 1138
rect 5038 1082 5050 1138
rect 4970 1048 5050 1082
rect 4970 992 4982 1048
rect 5038 992 5050 1048
rect 4970 958 5050 992
rect 4970 902 4982 958
rect 5038 902 5050 958
rect 4970 868 5050 902
rect 4970 812 4982 868
rect 5038 812 5050 868
rect 4970 800 5050 812
rect 5270 1318 5350 1340
rect 5270 1262 5282 1318
rect 5338 1262 5350 1318
rect 5270 1228 5350 1262
rect 5270 1172 5282 1228
rect 5338 1172 5350 1228
rect 5270 1138 5350 1172
rect 5270 1082 5282 1138
rect 5338 1082 5350 1138
rect 5270 1048 5350 1082
rect 5270 992 5282 1048
rect 5338 992 5350 1048
rect 5270 958 5350 992
rect 5270 902 5282 958
rect 5338 902 5350 958
rect 5270 868 5350 902
rect 5270 812 5282 868
rect 5338 812 5350 868
rect 5270 800 5350 812
rect 5570 1318 5650 1340
rect 5570 1262 5582 1318
rect 5638 1262 5650 1318
rect 5570 1228 5650 1262
rect 5570 1172 5582 1228
rect 5638 1172 5650 1228
rect 5570 1138 5650 1172
rect 5570 1082 5582 1138
rect 5638 1082 5650 1138
rect 5570 1048 5650 1082
rect 5570 992 5582 1048
rect 5638 992 5650 1048
rect 5570 958 5650 992
rect 5570 902 5582 958
rect 5638 902 5650 958
rect 5570 868 5650 902
rect 5570 812 5582 868
rect 5638 812 5650 868
rect 5570 800 5650 812
rect 5870 1318 5950 1340
rect 5870 1262 5882 1318
rect 5938 1262 5950 1318
rect 5870 1228 5950 1262
rect 5870 1172 5882 1228
rect 5938 1172 5950 1228
rect 5870 1138 5950 1172
rect 5870 1082 5882 1138
rect 5938 1082 5950 1138
rect 5870 1048 5950 1082
rect 5870 992 5882 1048
rect 5938 992 5950 1048
rect 5870 958 5950 992
rect 5870 902 5882 958
rect 5938 902 5950 958
rect 5870 868 5950 902
rect 5870 812 5882 868
rect 5938 812 5950 868
rect 5870 800 5950 812
rect 6170 1318 6250 1340
rect 6170 1262 6182 1318
rect 6238 1262 6250 1318
rect 6170 1228 6250 1262
rect 6170 1172 6182 1228
rect 6238 1172 6250 1228
rect 6170 1138 6250 1172
rect 6170 1082 6182 1138
rect 6238 1082 6250 1138
rect 6170 1048 6250 1082
rect 6170 992 6182 1048
rect 6238 992 6250 1048
rect 6170 958 6250 992
rect 6170 902 6182 958
rect 6238 902 6250 958
rect 6170 868 6250 902
rect 6170 812 6182 868
rect 6238 812 6250 868
rect 6170 800 6250 812
rect 490 390 550 800
rect 790 390 850 800
rect 1090 390 1150 800
rect 1390 390 1450 800
rect 1690 390 1750 800
rect 1990 390 2050 800
rect 2290 390 2350 800
rect 2590 390 2650 800
rect 2890 390 2950 800
rect 3490 390 3550 800
rect 3790 390 3850 800
rect 4090 390 4150 800
rect 4390 390 4450 800
rect 4690 390 4750 800
rect 4990 390 5050 800
rect 5290 390 5350 800
rect 5590 390 5650 800
rect 5890 390 5950 800
rect 6190 390 6250 800
rect 6570 2518 6650 2530
rect 6570 2462 6582 2518
rect 6638 2462 6650 2518
rect 6570 2428 6650 2462
rect 6570 2372 6582 2428
rect 6638 2372 6650 2428
rect -70 142 -58 198
rect -2 142 10 198
rect -70 108 10 142
rect -70 52 -58 108
rect -2 52 10 108
rect -70 -222 10 52
rect -70 -278 -58 -222
rect -2 -278 10 -222
rect -70 -312 10 -278
rect -70 -368 -58 -312
rect -2 -368 10 -312
rect 6570 198 6650 2372
rect 6570 142 6582 198
rect 6638 142 6650 198
rect 6570 108 6650 142
rect 6570 52 6582 108
rect 6638 52 6650 108
rect 6570 -222 6650 52
rect 6570 -278 6582 -222
rect 6638 -278 6650 -222
rect 6570 -312 6650 -278
rect 6570 -320 6582 -312
rect -70 -380 10 -368
rect 6460 -368 6582 -320
rect 6638 -368 6650 -312
rect 6460 -380 6650 -368
rect 6710 2428 6790 2440
rect 6710 2372 6722 2428
rect 6778 2372 6790 2428
rect 6710 2338 6790 2372
rect 6710 2282 6722 2338
rect 6778 2282 6790 2338
rect 6710 108 6790 2282
rect 6710 52 6722 108
rect 6778 52 6790 108
rect 6710 18 6790 52
rect 6710 -38 6722 18
rect 6778 -38 6790 18
rect 6710 -312 6790 -38
rect 6710 -368 6722 -312
rect 6778 -368 6790 -312
rect -210 -458 -198 -402
rect -142 -458 -130 -402
rect -210 -470 -130 -458
rect 6460 -590 6540 -380
rect 6710 -402 6790 -368
rect 6710 -458 6722 -402
rect 6778 -458 6790 -402
rect 6710 -590 6790 -458
rect 6447 -690 6557 -590
rect 6697 -690 6807 -590
<< via3 >>
rect 488 4978 552 5042
rect 788 4978 852 5042
rect 1088 4978 1152 5042
rect 1388 4978 1452 5042
rect 1688 4978 1752 5042
rect 1988 4978 2052 5042
rect 2288 4978 2352 5042
rect 2588 4978 2652 5042
rect 2888 4978 2952 5042
rect 3188 4978 3252 5042
rect 3488 4978 3552 5042
rect 3788 4978 3852 5042
rect 4088 4978 4152 5042
rect 4388 4978 4452 5042
rect 4688 4978 4752 5042
rect 4988 4978 5052 5042
rect 5288 4978 5352 5042
rect 5588 4978 5652 5042
rect 5888 4978 5952 5042
rect 6188 4978 6252 5042
<< metal4 >>
rect -493 5042 6897 5060
rect -493 4978 488 5042
rect 552 4978 788 5042
rect 852 4978 1088 5042
rect 1152 4978 1388 5042
rect 1452 4978 1688 5042
rect 1752 4978 1988 5042
rect 2052 4978 2288 5042
rect 2352 4978 2588 5042
rect 2652 4978 2888 5042
rect 2952 4978 3188 5042
rect 3252 4978 3488 5042
rect 3552 4978 3788 5042
rect 3852 4978 4088 5042
rect 4152 4978 4388 5042
rect 4452 4978 4688 5042
rect 4752 4978 4988 5042
rect 5052 4978 5288 5042
rect 5352 4978 5588 5042
rect 5652 4978 5888 5042
rect 5952 4978 6188 5042
rect 6252 4978 6897 5042
rect -493 4960 6897 4978
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_0
timestamp 1757161594
transform 0 1 1648 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_1
timestamp 1757161594
transform 0 1 1348 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_2
timestamp 1757161594
transform 0 1 448 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_3
timestamp 1757161594
transform 0 1 148 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_4
timestamp 1757161594
transform 0 1 1048 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_5
timestamp 1757161594
transform 0 1 748 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_6
timestamp 1757161594
transform 0 1 2848 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_7
timestamp 1757161594
transform 0 1 3148 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_8
timestamp 1757161594
transform 0 1 2248 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_9
timestamp 1757161594
transform 0 1 2548 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_10
timestamp 1757161594
transform 0 1 1948 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_11
timestamp 1757161594
transform 0 1 3448 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_12
timestamp 1757161594
transform 0 1 4648 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_13
timestamp 1757161594
transform 0 1 4948 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_14
timestamp 1757161594
transform 0 1 4048 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_15
timestamp 1757161594
transform 0 1 4348 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_16
timestamp 1757161594
transform 0 1 3748 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_17
timestamp 1757161594
transform 0 1 5248 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_18
timestamp 1757161594
transform 0 1 6448 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_19
timestamp 1757161594
transform 0 1 5848 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_20
timestamp 1757161594
transform 0 1 6148 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_21
timestamp 1757161594
transform 0 1 5548 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_22
timestamp 1757161594
transform 0 1 1648 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_23
timestamp 1757161594
transform 0 1 1348 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_24
timestamp 1757161594
transform 0 1 1048 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_25
timestamp 1757161594
transform 0 1 748 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_26
timestamp 1757161594
transform 0 1 448 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_28
timestamp 1757161594
transform 0 1 1948 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_29
timestamp 1757161594
transform 0 1 2248 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_30
timestamp 1757161594
transform 0 1 2548 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_31
timestamp 1757161594
transform 0 1 2848 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_32
timestamp 1757161594
transform 0 1 3148 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_33
timestamp 1757161594
transform 0 1 3448 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_34
timestamp 1757161594
transform 0 1 3748 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_35
timestamp 1757161594
transform 0 1 4048 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_36
timestamp 1757161594
transform 0 1 4348 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_37
timestamp 1757161594
transform 0 1 4648 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_38
timestamp 1757161594
transform 0 1 4948 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_39
timestamp 1757161594
transform 0 1 5248 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_40
timestamp 1757161594
transform 0 1 5548 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_41
timestamp 1757161594
transform 0 1 5848 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_42
timestamp 1757161594
transform 0 1 6148 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_43
timestamp 1757161594
transform 0 1 6448 1 0 -186
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSMGKB  sky130_fd_pr__pfet_01v8_lvt_RSMGKB_44
timestamp 1757161594
transform 0 1 148 1 0 4694
box -144 -148 144 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_0
timestamp 1757161594
transform 0 1 2848 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_1
timestamp 1757161594
transform 0 1 1648 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_2
timestamp 1757161594
transform 0 1 1948 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_3
timestamp 1757161594
transform 0 1 2248 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_4
timestamp 1757161594
transform 0 1 2548 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_5
timestamp 1757161594
transform 0 1 1348 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_6
timestamp 1757161594
transform 0 1 1048 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_7
timestamp 1757161594
transform 0 1 748 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_8
timestamp 1757161594
transform 0 1 448 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_9
timestamp 1757161594
transform 0 1 448 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_10
timestamp 1757161594
transform 0 1 4648 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_11
timestamp 1757161594
transform 0 1 4948 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_12
timestamp 1757161594
transform 0 1 5248 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_13
timestamp 1757161594
transform 0 1 5548 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_14
timestamp 1757161594
transform 0 1 5848 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_15
timestamp 1757161594
transform 0 1 3148 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_16
timestamp 1757161594
transform 0 1 3448 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_17
timestamp 1757161594
transform 0 1 3748 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_18
timestamp 1757161594
transform 0 1 4048 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_19
timestamp 1757161594
transform 0 1 4348 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_20
timestamp 1757161594
transform 0 1 6148 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_21
timestamp 1757161594
transform 0 1 6448 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_22
timestamp 1757161594
transform 0 1 148 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_23
timestamp 1757161594
transform 0 1 148 1 0 1094
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_44
timestamp 1757161594
transform 0 1 1648 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_45
timestamp 1757161594
transform 0 1 1348 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_46
timestamp 1757161594
transform 0 1 1048 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_47
timestamp 1757161594
transform 0 1 748 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_50
timestamp 1757161594
transform 0 1 3148 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_51
timestamp 1757161594
transform 0 1 2848 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_52
timestamp 1757161594
transform 0 1 2548 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_53
timestamp 1757161594
transform 0 1 2248 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_54
timestamp 1757161594
transform 0 1 1948 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_55
timestamp 1757161594
transform 0 1 4948 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_56
timestamp 1757161594
transform 0 1 4648 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_57
timestamp 1757161594
transform 0 1 4348 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_58
timestamp 1757161594
transform 0 1 4048 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_59
timestamp 1757161594
transform 0 1 3748 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_60
timestamp 1757161594
transform 0 1 3448 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_61
timestamp 1757161594
transform 0 1 6448 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_62
timestamp 1757161594
transform 0 1 6148 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_63
timestamp 1757161594
transform 0 1 5848 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_64
timestamp 1757161594
transform 0 1 5548 1 0 3414
box -1094 -148 1094 114
use sky130_fd_pr__pfet_01v8_lvt_RSW4TG  sky130_fd_pr__pfet_01v8_lvt_RSW4TG_65
timestamp 1757161594
transform 0 1 5248 1 0 3414
box -1094 -148 1094 114
<< labels >>
flabel metal4 s -493 4960 -413 5060 0 FreeSans 782 180 0 0 Vbin
port 0 nsew
<< end >>
