magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -343 5257 9003 5343
rect -343 60 -257 5257
rect -343 -90 -24 60
rect 4064 -60 4156 80
rect -343 -5157 -257 -90
rect 8917 -5157 9003 5257
rect -343 -5243 9003 -5157
<< psubdiff >>
rect -317 5283 -243 5317
rect -209 5283 -175 5317
rect -141 5283 -107 5317
rect -73 5283 -39 5317
rect -5 5283 29 5317
rect 63 5283 97 5317
rect 131 5283 165 5317
rect 199 5283 233 5317
rect 267 5283 301 5317
rect 335 5283 369 5317
rect 403 5283 437 5317
rect 471 5283 505 5317
rect 539 5283 573 5317
rect 607 5283 641 5317
rect 675 5283 709 5317
rect 743 5283 777 5317
rect 811 5283 845 5317
rect 879 5283 913 5317
rect 947 5283 981 5317
rect 1015 5283 1049 5317
rect 1083 5283 1117 5317
rect 1151 5283 1185 5317
rect 1219 5283 1253 5317
rect 1287 5283 1321 5317
rect 1355 5283 1389 5317
rect 1423 5283 1457 5317
rect 1491 5283 1525 5317
rect 1559 5283 1593 5317
rect 1627 5283 1661 5317
rect 1695 5283 1729 5317
rect 1763 5283 1797 5317
rect 1831 5283 1865 5317
rect 1899 5283 1933 5317
rect 1967 5283 2001 5317
rect 2035 5283 2069 5317
rect 2103 5283 2137 5317
rect 2171 5283 2205 5317
rect 2239 5283 2273 5317
rect 2307 5283 2341 5317
rect 2375 5283 2409 5317
rect 2443 5283 2477 5317
rect 2511 5283 2545 5317
rect 2579 5283 2613 5317
rect 2647 5283 2681 5317
rect 2715 5283 2749 5317
rect 2783 5283 2817 5317
rect 2851 5283 2885 5317
rect 2919 5283 2953 5317
rect 2987 5283 3021 5317
rect 3055 5283 3089 5317
rect 3123 5283 3157 5317
rect 3191 5283 3225 5317
rect 3259 5283 3293 5317
rect 3327 5283 3361 5317
rect 3395 5283 3429 5317
rect 3463 5283 3497 5317
rect 3531 5283 3565 5317
rect 3599 5283 3633 5317
rect 3667 5283 3701 5317
rect 3735 5283 3769 5317
rect 3803 5283 3837 5317
rect 3871 5283 3905 5317
rect 3939 5283 3973 5317
rect 4007 5283 4041 5317
rect 4075 5283 4109 5317
rect 4143 5283 4177 5317
rect 4211 5283 4245 5317
rect 4279 5283 4313 5317
rect 4347 5283 4381 5317
rect 4415 5283 4449 5317
rect 4483 5283 4517 5317
rect 4551 5283 4585 5317
rect 4619 5283 4653 5317
rect 4687 5283 4721 5317
rect 4755 5283 4789 5317
rect 4823 5283 4857 5317
rect 4891 5283 4925 5317
rect 4959 5283 4993 5317
rect 5027 5283 5061 5317
rect 5095 5283 5129 5317
rect 5163 5283 5197 5317
rect 5231 5283 5265 5317
rect 5299 5283 5333 5317
rect 5367 5283 5401 5317
rect 5435 5283 5469 5317
rect 5503 5283 5537 5317
rect 5571 5283 5605 5317
rect 5639 5283 5673 5317
rect 5707 5283 5741 5317
rect 5775 5283 5809 5317
rect 5843 5283 5877 5317
rect 5911 5283 5945 5317
rect 5979 5283 6013 5317
rect 6047 5283 6081 5317
rect 6115 5283 6149 5317
rect 6183 5283 6217 5317
rect 6251 5283 6285 5317
rect 6319 5283 6353 5317
rect 6387 5283 6421 5317
rect 6455 5283 6489 5317
rect 6523 5283 6557 5317
rect 6591 5283 6625 5317
rect 6659 5283 6693 5317
rect 6727 5283 6761 5317
rect 6795 5283 6829 5317
rect 6863 5283 6897 5317
rect 6931 5283 6965 5317
rect 6999 5283 7033 5317
rect 7067 5283 7101 5317
rect 7135 5283 7169 5317
rect 7203 5283 7237 5317
rect 7271 5283 7305 5317
rect 7339 5283 7373 5317
rect 7407 5283 7441 5317
rect 7475 5283 7509 5317
rect 7543 5283 7577 5317
rect 7611 5283 7645 5317
rect 7679 5283 7713 5317
rect 7747 5283 7781 5317
rect 7815 5283 7849 5317
rect 7883 5283 7917 5317
rect 7951 5283 7985 5317
rect 8019 5283 8053 5317
rect 8087 5283 8121 5317
rect 8155 5283 8189 5317
rect 8223 5283 8257 5317
rect 8291 5283 8325 5317
rect 8359 5283 8393 5317
rect 8427 5283 8461 5317
rect 8495 5283 8529 5317
rect 8563 5283 8597 5317
rect 8631 5283 8665 5317
rect 8699 5283 8733 5317
rect 8767 5283 8801 5317
rect 8835 5283 8869 5317
rect 8903 5283 8977 5317
rect -317 5235 -283 5283
rect -317 5167 -283 5201
rect -317 5099 -283 5133
rect -317 5031 -283 5065
rect -317 4963 -283 4997
rect -317 4895 -283 4929
rect -317 4827 -283 4861
rect -317 4759 -283 4793
rect -317 4691 -283 4725
rect -317 4623 -283 4657
rect -317 4555 -283 4589
rect -317 4487 -283 4521
rect -317 4419 -283 4453
rect -317 4351 -283 4385
rect -317 4283 -283 4317
rect -317 4215 -283 4249
rect -317 4147 -283 4181
rect -317 4079 -283 4113
rect -317 4011 -283 4045
rect -317 3943 -283 3977
rect -317 3875 -283 3909
rect -317 3807 -283 3841
rect -317 3739 -283 3773
rect -317 3671 -283 3705
rect -317 3603 -283 3637
rect -317 3535 -283 3569
rect -317 3467 -283 3501
rect -317 3399 -283 3433
rect -317 3331 -283 3365
rect -317 3263 -283 3297
rect -317 3195 -283 3229
rect -317 3127 -283 3161
rect -317 3059 -283 3093
rect -317 2991 -283 3025
rect -317 2923 -283 2957
rect -317 2855 -283 2889
rect -317 2787 -283 2821
rect -317 2719 -283 2753
rect -317 2651 -283 2685
rect -317 2583 -283 2617
rect -317 2515 -283 2549
rect -317 2447 -283 2481
rect -317 2379 -283 2413
rect -317 2311 -283 2345
rect -317 2243 -283 2277
rect -317 2175 -283 2209
rect -317 2107 -283 2141
rect -317 2039 -283 2073
rect -317 1971 -283 2005
rect -317 1903 -283 1937
rect -317 1835 -283 1869
rect -317 1767 -283 1801
rect -317 1699 -283 1733
rect -317 1631 -283 1665
rect -317 1563 -283 1597
rect -317 1495 -283 1529
rect -317 1427 -283 1461
rect -317 1359 -283 1393
rect -317 1291 -283 1325
rect -317 1223 -283 1257
rect -317 1155 -283 1189
rect -317 1087 -283 1121
rect -317 1019 -283 1053
rect -317 951 -283 985
rect -317 883 -283 917
rect -317 815 -283 849
rect -317 747 -283 781
rect -317 679 -283 713
rect -317 611 -283 645
rect -317 543 -283 577
rect -317 475 -283 509
rect -317 407 -283 441
rect -317 339 -283 373
rect -317 271 -283 305
rect -317 203 -283 237
rect -317 135 -283 169
rect -317 67 -283 101
rect 8943 5235 8977 5283
rect 8943 5167 8977 5201
rect 8943 5099 8977 5133
rect 8943 5031 8977 5065
rect 8943 4963 8977 4997
rect 8943 4895 8977 4929
rect 8943 4827 8977 4861
rect 8943 4759 8977 4793
rect 8943 4691 8977 4725
rect 8943 4623 8977 4657
rect 8943 4555 8977 4589
rect 8943 4487 8977 4521
rect 8943 4419 8977 4453
rect 8943 4351 8977 4385
rect 8943 4283 8977 4317
rect 8943 4215 8977 4249
rect 8943 4147 8977 4181
rect 8943 4079 8977 4113
rect 8943 4011 8977 4045
rect 8943 3943 8977 3977
rect 8943 3875 8977 3909
rect 8943 3807 8977 3841
rect 8943 3739 8977 3773
rect 8943 3671 8977 3705
rect 8943 3603 8977 3637
rect 8943 3535 8977 3569
rect 8943 3467 8977 3501
rect 8943 3399 8977 3433
rect 8943 3331 8977 3365
rect 8943 3263 8977 3297
rect 8943 3195 8977 3229
rect 8943 3127 8977 3161
rect 8943 3059 8977 3093
rect 8943 2991 8977 3025
rect 8943 2923 8977 2957
rect 8943 2855 8977 2889
rect 8943 2787 8977 2821
rect 8943 2719 8977 2753
rect 8943 2651 8977 2685
rect 8943 2583 8977 2617
rect 8943 2515 8977 2549
rect 8943 2447 8977 2481
rect 8943 2379 8977 2413
rect 8943 2311 8977 2345
rect 8943 2243 8977 2277
rect 8943 2175 8977 2209
rect 8943 2107 8977 2141
rect 8943 2039 8977 2073
rect 8943 1971 8977 2005
rect 8943 1903 8977 1937
rect 8943 1835 8977 1869
rect 8943 1767 8977 1801
rect 8943 1699 8977 1733
rect 8943 1631 8977 1665
rect 8943 1563 8977 1597
rect 8943 1495 8977 1529
rect 8943 1427 8977 1461
rect 8943 1359 8977 1393
rect 8943 1291 8977 1325
rect 8943 1223 8977 1257
rect 8943 1155 8977 1189
rect 8943 1087 8977 1121
rect 8943 1019 8977 1053
rect 8943 951 8977 985
rect 8943 883 8977 917
rect 8943 815 8977 849
rect 8943 747 8977 781
rect 8943 679 8977 713
rect 8943 611 8977 645
rect 8943 543 8977 577
rect 8943 475 8977 509
rect 8943 407 8977 441
rect 8943 339 8977 373
rect 8943 271 8977 305
rect 8943 203 8977 237
rect 8943 135 8977 169
rect 8943 67 8977 101
rect -317 -1 -283 33
rect -317 -69 -283 -35
rect -100 2 -50 34
rect -100 -32 -92 2
rect -58 -32 -50 2
rect -100 -64 -50 -32
rect 4090 27 4130 54
rect 4090 -7 4093 27
rect 4127 -7 4130 27
rect 4090 -34 4130 -7
rect 8943 -1 8977 33
rect -317 -137 -283 -103
rect -317 -205 -283 -171
rect -317 -273 -283 -239
rect -317 -341 -283 -307
rect -317 -409 -283 -375
rect -317 -477 -283 -443
rect -317 -545 -283 -511
rect -317 -613 -283 -579
rect -317 -681 -283 -647
rect -317 -749 -283 -715
rect -317 -817 -283 -783
rect -317 -885 -283 -851
rect -317 -953 -283 -919
rect -317 -1021 -283 -987
rect -317 -1089 -283 -1055
rect -317 -1157 -283 -1123
rect -317 -1225 -283 -1191
rect -317 -1293 -283 -1259
rect -317 -1361 -283 -1327
rect -317 -1429 -283 -1395
rect -317 -1497 -283 -1463
rect -317 -1565 -283 -1531
rect -317 -1633 -283 -1599
rect -317 -1701 -283 -1667
rect -317 -1769 -283 -1735
rect -317 -1837 -283 -1803
rect -317 -1905 -283 -1871
rect -317 -1973 -283 -1939
rect -317 -2041 -283 -2007
rect -317 -2109 -283 -2075
rect -317 -2177 -283 -2143
rect -317 -2245 -283 -2211
rect -317 -2313 -283 -2279
rect -317 -2381 -283 -2347
rect -317 -2449 -283 -2415
rect -317 -2517 -283 -2483
rect -317 -2585 -283 -2551
rect -317 -2653 -283 -2619
rect -317 -2721 -283 -2687
rect -317 -2789 -283 -2755
rect -317 -2857 -283 -2823
rect -317 -2925 -283 -2891
rect -317 -2993 -283 -2959
rect -317 -3061 -283 -3027
rect -317 -3129 -283 -3095
rect -317 -3197 -283 -3163
rect -317 -3265 -283 -3231
rect -317 -3333 -283 -3299
rect -317 -3401 -283 -3367
rect -317 -3469 -283 -3435
rect -317 -3537 -283 -3503
rect -317 -3605 -283 -3571
rect -317 -3673 -283 -3639
rect -317 -3741 -283 -3707
rect -317 -3809 -283 -3775
rect -317 -3877 -283 -3843
rect -317 -3945 -283 -3911
rect -317 -4013 -283 -3979
rect -317 -4081 -283 -4047
rect -317 -4149 -283 -4115
rect -317 -4217 -283 -4183
rect -317 -4285 -283 -4251
rect -317 -4353 -283 -4319
rect -317 -4421 -283 -4387
rect -317 -4489 -283 -4455
rect -317 -4557 -283 -4523
rect -317 -4625 -283 -4591
rect -317 -4693 -283 -4659
rect -317 -4761 -283 -4727
rect -317 -4829 -283 -4795
rect -317 -4897 -283 -4863
rect -317 -4965 -283 -4931
rect -317 -5033 -283 -4999
rect -317 -5101 -283 -5067
rect -317 -5183 -283 -5135
rect 8943 -69 8977 -35
rect 8943 -137 8977 -103
rect 8943 -205 8977 -171
rect 8943 -273 8977 -239
rect 8943 -341 8977 -307
rect 8943 -409 8977 -375
rect 8943 -477 8977 -443
rect 8943 -545 8977 -511
rect 8943 -613 8977 -579
rect 8943 -681 8977 -647
rect 8943 -749 8977 -715
rect 8943 -817 8977 -783
rect 8943 -885 8977 -851
rect 8943 -953 8977 -919
rect 8943 -1021 8977 -987
rect 8943 -1089 8977 -1055
rect 8943 -1157 8977 -1123
rect 8943 -1225 8977 -1191
rect 8943 -1293 8977 -1259
rect 8943 -1361 8977 -1327
rect 8943 -1429 8977 -1395
rect 8943 -1497 8977 -1463
rect 8943 -1565 8977 -1531
rect 8943 -1633 8977 -1599
rect 8943 -1701 8977 -1667
rect 8943 -1769 8977 -1735
rect 8943 -1837 8977 -1803
rect 8943 -1905 8977 -1871
rect 8943 -1973 8977 -1939
rect 8943 -2041 8977 -2007
rect 8943 -2109 8977 -2075
rect 8943 -2177 8977 -2143
rect 8943 -2245 8977 -2211
rect 8943 -2313 8977 -2279
rect 8943 -2381 8977 -2347
rect 8943 -2449 8977 -2415
rect 8943 -2517 8977 -2483
rect 8943 -2585 8977 -2551
rect 8943 -2653 8977 -2619
rect 8943 -2721 8977 -2687
rect 8943 -2789 8977 -2755
rect 8943 -2857 8977 -2823
rect 8943 -2925 8977 -2891
rect 8943 -2993 8977 -2959
rect 8943 -3061 8977 -3027
rect 8943 -3129 8977 -3095
rect 8943 -3197 8977 -3163
rect 8943 -3265 8977 -3231
rect 8943 -3333 8977 -3299
rect 8943 -3401 8977 -3367
rect 8943 -3469 8977 -3435
rect 8943 -3537 8977 -3503
rect 8943 -3605 8977 -3571
rect 8943 -3673 8977 -3639
rect 8943 -3741 8977 -3707
rect 8943 -3809 8977 -3775
rect 8943 -3877 8977 -3843
rect 8943 -3945 8977 -3911
rect 8943 -4013 8977 -3979
rect 8943 -4081 8977 -4047
rect 8943 -4149 8977 -4115
rect 8943 -4217 8977 -4183
rect 8943 -4285 8977 -4251
rect 8943 -4353 8977 -4319
rect 8943 -4421 8977 -4387
rect 8943 -4489 8977 -4455
rect 8943 -4557 8977 -4523
rect 8943 -4625 8977 -4591
rect 8943 -4693 8977 -4659
rect 8943 -4761 8977 -4727
rect 8943 -4829 8977 -4795
rect 8943 -4897 8977 -4863
rect 8943 -4965 8977 -4931
rect 8943 -5033 8977 -4999
rect 8943 -5101 8977 -5067
rect 8943 -5183 8977 -5135
rect -317 -5217 -243 -5183
rect -209 -5217 -175 -5183
rect -141 -5217 -107 -5183
rect -73 -5217 -39 -5183
rect -5 -5217 29 -5183
rect 63 -5217 97 -5183
rect 131 -5217 165 -5183
rect 199 -5217 233 -5183
rect 267 -5217 301 -5183
rect 335 -5217 369 -5183
rect 403 -5217 437 -5183
rect 471 -5217 505 -5183
rect 539 -5217 573 -5183
rect 607 -5217 641 -5183
rect 675 -5217 709 -5183
rect 743 -5217 777 -5183
rect 811 -5217 845 -5183
rect 879 -5217 913 -5183
rect 947 -5217 981 -5183
rect 1015 -5217 1049 -5183
rect 1083 -5217 1117 -5183
rect 1151 -5217 1185 -5183
rect 1219 -5217 1253 -5183
rect 1287 -5217 1321 -5183
rect 1355 -5217 1389 -5183
rect 1423 -5217 1457 -5183
rect 1491 -5217 1525 -5183
rect 1559 -5217 1593 -5183
rect 1627 -5217 1661 -5183
rect 1695 -5217 1729 -5183
rect 1763 -5217 1797 -5183
rect 1831 -5217 1865 -5183
rect 1899 -5217 1933 -5183
rect 1967 -5217 2001 -5183
rect 2035 -5217 2069 -5183
rect 2103 -5217 2137 -5183
rect 2171 -5217 2205 -5183
rect 2239 -5217 2273 -5183
rect 2307 -5217 2341 -5183
rect 2375 -5217 2409 -5183
rect 2443 -5217 2477 -5183
rect 2511 -5217 2545 -5183
rect 2579 -5217 2613 -5183
rect 2647 -5217 2681 -5183
rect 2715 -5217 2749 -5183
rect 2783 -5217 2817 -5183
rect 2851 -5217 2885 -5183
rect 2919 -5217 2953 -5183
rect 2987 -5217 3021 -5183
rect 3055 -5217 3089 -5183
rect 3123 -5217 3157 -5183
rect 3191 -5217 3225 -5183
rect 3259 -5217 3293 -5183
rect 3327 -5217 3361 -5183
rect 3395 -5217 3429 -5183
rect 3463 -5217 3497 -5183
rect 3531 -5217 3565 -5183
rect 3599 -5217 3633 -5183
rect 3667 -5217 3701 -5183
rect 3735 -5217 3769 -5183
rect 3803 -5217 3837 -5183
rect 3871 -5217 3905 -5183
rect 3939 -5217 3973 -5183
rect 4007 -5217 4041 -5183
rect 4075 -5217 4109 -5183
rect 4143 -5217 4177 -5183
rect 4211 -5217 4245 -5183
rect 4279 -5217 4313 -5183
rect 4347 -5217 4381 -5183
rect 4415 -5217 4449 -5183
rect 4483 -5217 4517 -5183
rect 4551 -5217 4585 -5183
rect 4619 -5217 4653 -5183
rect 4687 -5217 4721 -5183
rect 4755 -5217 4789 -5183
rect 4823 -5217 4857 -5183
rect 4891 -5217 4925 -5183
rect 4959 -5217 4993 -5183
rect 5027 -5217 5061 -5183
rect 5095 -5217 5129 -5183
rect 5163 -5217 5197 -5183
rect 5231 -5217 5265 -5183
rect 5299 -5217 5333 -5183
rect 5367 -5217 5401 -5183
rect 5435 -5217 5469 -5183
rect 5503 -5217 5537 -5183
rect 5571 -5217 5605 -5183
rect 5639 -5217 5673 -5183
rect 5707 -5217 5741 -5183
rect 5775 -5217 5809 -5183
rect 5843 -5217 5877 -5183
rect 5911 -5217 5945 -5183
rect 5979 -5217 6013 -5183
rect 6047 -5217 6081 -5183
rect 6115 -5217 6149 -5183
rect 6183 -5217 6217 -5183
rect 6251 -5217 6285 -5183
rect 6319 -5217 6353 -5183
rect 6387 -5217 6421 -5183
rect 6455 -5217 6489 -5183
rect 6523 -5217 6557 -5183
rect 6591 -5217 6625 -5183
rect 6659 -5217 6693 -5183
rect 6727 -5217 6761 -5183
rect 6795 -5217 6829 -5183
rect 6863 -5217 6897 -5183
rect 6931 -5217 6965 -5183
rect 6999 -5217 7033 -5183
rect 7067 -5217 7101 -5183
rect 7135 -5217 7169 -5183
rect 7203 -5217 7237 -5183
rect 7271 -5217 7305 -5183
rect 7339 -5217 7373 -5183
rect 7407 -5217 7441 -5183
rect 7475 -5217 7509 -5183
rect 7543 -5217 7577 -5183
rect 7611 -5217 7645 -5183
rect 7679 -5217 7713 -5183
rect 7747 -5217 7781 -5183
rect 7815 -5217 7849 -5183
rect 7883 -5217 7917 -5183
rect 7951 -5217 7985 -5183
rect 8019 -5217 8053 -5183
rect 8087 -5217 8121 -5183
rect 8155 -5217 8189 -5183
rect 8223 -5217 8257 -5183
rect 8291 -5217 8325 -5183
rect 8359 -5217 8393 -5183
rect 8427 -5217 8461 -5183
rect 8495 -5217 8529 -5183
rect 8563 -5217 8597 -5183
rect 8631 -5217 8665 -5183
rect 8699 -5217 8733 -5183
rect 8767 -5217 8801 -5183
rect 8835 -5217 8869 -5183
rect 8903 -5217 8977 -5183
<< psubdiffcont >>
rect -243 5283 -209 5317
rect -175 5283 -141 5317
rect -107 5283 -73 5317
rect -39 5283 -5 5317
rect 29 5283 63 5317
rect 97 5283 131 5317
rect 165 5283 199 5317
rect 233 5283 267 5317
rect 301 5283 335 5317
rect 369 5283 403 5317
rect 437 5283 471 5317
rect 505 5283 539 5317
rect 573 5283 607 5317
rect 641 5283 675 5317
rect 709 5283 743 5317
rect 777 5283 811 5317
rect 845 5283 879 5317
rect 913 5283 947 5317
rect 981 5283 1015 5317
rect 1049 5283 1083 5317
rect 1117 5283 1151 5317
rect 1185 5283 1219 5317
rect 1253 5283 1287 5317
rect 1321 5283 1355 5317
rect 1389 5283 1423 5317
rect 1457 5283 1491 5317
rect 1525 5283 1559 5317
rect 1593 5283 1627 5317
rect 1661 5283 1695 5317
rect 1729 5283 1763 5317
rect 1797 5283 1831 5317
rect 1865 5283 1899 5317
rect 1933 5283 1967 5317
rect 2001 5283 2035 5317
rect 2069 5283 2103 5317
rect 2137 5283 2171 5317
rect 2205 5283 2239 5317
rect 2273 5283 2307 5317
rect 2341 5283 2375 5317
rect 2409 5283 2443 5317
rect 2477 5283 2511 5317
rect 2545 5283 2579 5317
rect 2613 5283 2647 5317
rect 2681 5283 2715 5317
rect 2749 5283 2783 5317
rect 2817 5283 2851 5317
rect 2885 5283 2919 5317
rect 2953 5283 2987 5317
rect 3021 5283 3055 5317
rect 3089 5283 3123 5317
rect 3157 5283 3191 5317
rect 3225 5283 3259 5317
rect 3293 5283 3327 5317
rect 3361 5283 3395 5317
rect 3429 5283 3463 5317
rect 3497 5283 3531 5317
rect 3565 5283 3599 5317
rect 3633 5283 3667 5317
rect 3701 5283 3735 5317
rect 3769 5283 3803 5317
rect 3837 5283 3871 5317
rect 3905 5283 3939 5317
rect 3973 5283 4007 5317
rect 4041 5283 4075 5317
rect 4109 5283 4143 5317
rect 4177 5283 4211 5317
rect 4245 5283 4279 5317
rect 4313 5283 4347 5317
rect 4381 5283 4415 5317
rect 4449 5283 4483 5317
rect 4517 5283 4551 5317
rect 4585 5283 4619 5317
rect 4653 5283 4687 5317
rect 4721 5283 4755 5317
rect 4789 5283 4823 5317
rect 4857 5283 4891 5317
rect 4925 5283 4959 5317
rect 4993 5283 5027 5317
rect 5061 5283 5095 5317
rect 5129 5283 5163 5317
rect 5197 5283 5231 5317
rect 5265 5283 5299 5317
rect 5333 5283 5367 5317
rect 5401 5283 5435 5317
rect 5469 5283 5503 5317
rect 5537 5283 5571 5317
rect 5605 5283 5639 5317
rect 5673 5283 5707 5317
rect 5741 5283 5775 5317
rect 5809 5283 5843 5317
rect 5877 5283 5911 5317
rect 5945 5283 5979 5317
rect 6013 5283 6047 5317
rect 6081 5283 6115 5317
rect 6149 5283 6183 5317
rect 6217 5283 6251 5317
rect 6285 5283 6319 5317
rect 6353 5283 6387 5317
rect 6421 5283 6455 5317
rect 6489 5283 6523 5317
rect 6557 5283 6591 5317
rect 6625 5283 6659 5317
rect 6693 5283 6727 5317
rect 6761 5283 6795 5317
rect 6829 5283 6863 5317
rect 6897 5283 6931 5317
rect 6965 5283 6999 5317
rect 7033 5283 7067 5317
rect 7101 5283 7135 5317
rect 7169 5283 7203 5317
rect 7237 5283 7271 5317
rect 7305 5283 7339 5317
rect 7373 5283 7407 5317
rect 7441 5283 7475 5317
rect 7509 5283 7543 5317
rect 7577 5283 7611 5317
rect 7645 5283 7679 5317
rect 7713 5283 7747 5317
rect 7781 5283 7815 5317
rect 7849 5283 7883 5317
rect 7917 5283 7951 5317
rect 7985 5283 8019 5317
rect 8053 5283 8087 5317
rect 8121 5283 8155 5317
rect 8189 5283 8223 5317
rect 8257 5283 8291 5317
rect 8325 5283 8359 5317
rect 8393 5283 8427 5317
rect 8461 5283 8495 5317
rect 8529 5283 8563 5317
rect 8597 5283 8631 5317
rect 8665 5283 8699 5317
rect 8733 5283 8767 5317
rect 8801 5283 8835 5317
rect 8869 5283 8903 5317
rect -317 5201 -283 5235
rect -317 5133 -283 5167
rect -317 5065 -283 5099
rect -317 4997 -283 5031
rect -317 4929 -283 4963
rect -317 4861 -283 4895
rect -317 4793 -283 4827
rect -317 4725 -283 4759
rect -317 4657 -283 4691
rect -317 4589 -283 4623
rect -317 4521 -283 4555
rect -317 4453 -283 4487
rect -317 4385 -283 4419
rect -317 4317 -283 4351
rect -317 4249 -283 4283
rect -317 4181 -283 4215
rect -317 4113 -283 4147
rect -317 4045 -283 4079
rect -317 3977 -283 4011
rect -317 3909 -283 3943
rect -317 3841 -283 3875
rect -317 3773 -283 3807
rect -317 3705 -283 3739
rect -317 3637 -283 3671
rect -317 3569 -283 3603
rect -317 3501 -283 3535
rect -317 3433 -283 3467
rect -317 3365 -283 3399
rect -317 3297 -283 3331
rect -317 3229 -283 3263
rect -317 3161 -283 3195
rect -317 3093 -283 3127
rect -317 3025 -283 3059
rect -317 2957 -283 2991
rect -317 2889 -283 2923
rect -317 2821 -283 2855
rect -317 2753 -283 2787
rect -317 2685 -283 2719
rect -317 2617 -283 2651
rect -317 2549 -283 2583
rect -317 2481 -283 2515
rect -317 2413 -283 2447
rect -317 2345 -283 2379
rect -317 2277 -283 2311
rect -317 2209 -283 2243
rect -317 2141 -283 2175
rect -317 2073 -283 2107
rect -317 2005 -283 2039
rect -317 1937 -283 1971
rect -317 1869 -283 1903
rect -317 1801 -283 1835
rect -317 1733 -283 1767
rect -317 1665 -283 1699
rect -317 1597 -283 1631
rect -317 1529 -283 1563
rect -317 1461 -283 1495
rect -317 1393 -283 1427
rect -317 1325 -283 1359
rect -317 1257 -283 1291
rect -317 1189 -283 1223
rect -317 1121 -283 1155
rect -317 1053 -283 1087
rect -317 985 -283 1019
rect -317 917 -283 951
rect -317 849 -283 883
rect -317 781 -283 815
rect -317 713 -283 747
rect -317 645 -283 679
rect -317 577 -283 611
rect -317 509 -283 543
rect -317 441 -283 475
rect -317 373 -283 407
rect -317 305 -283 339
rect -317 237 -283 271
rect -317 169 -283 203
rect -317 101 -283 135
rect -317 33 -283 67
rect 8943 5201 8977 5235
rect 8943 5133 8977 5167
rect 8943 5065 8977 5099
rect 8943 4997 8977 5031
rect 8943 4929 8977 4963
rect 8943 4861 8977 4895
rect 8943 4793 8977 4827
rect 8943 4725 8977 4759
rect 8943 4657 8977 4691
rect 8943 4589 8977 4623
rect 8943 4521 8977 4555
rect 8943 4453 8977 4487
rect 8943 4385 8977 4419
rect 8943 4317 8977 4351
rect 8943 4249 8977 4283
rect 8943 4181 8977 4215
rect 8943 4113 8977 4147
rect 8943 4045 8977 4079
rect 8943 3977 8977 4011
rect 8943 3909 8977 3943
rect 8943 3841 8977 3875
rect 8943 3773 8977 3807
rect 8943 3705 8977 3739
rect 8943 3637 8977 3671
rect 8943 3569 8977 3603
rect 8943 3501 8977 3535
rect 8943 3433 8977 3467
rect 8943 3365 8977 3399
rect 8943 3297 8977 3331
rect 8943 3229 8977 3263
rect 8943 3161 8977 3195
rect 8943 3093 8977 3127
rect 8943 3025 8977 3059
rect 8943 2957 8977 2991
rect 8943 2889 8977 2923
rect 8943 2821 8977 2855
rect 8943 2753 8977 2787
rect 8943 2685 8977 2719
rect 8943 2617 8977 2651
rect 8943 2549 8977 2583
rect 8943 2481 8977 2515
rect 8943 2413 8977 2447
rect 8943 2345 8977 2379
rect 8943 2277 8977 2311
rect 8943 2209 8977 2243
rect 8943 2141 8977 2175
rect 8943 2073 8977 2107
rect 8943 2005 8977 2039
rect 8943 1937 8977 1971
rect 8943 1869 8977 1903
rect 8943 1801 8977 1835
rect 8943 1733 8977 1767
rect 8943 1665 8977 1699
rect 8943 1597 8977 1631
rect 8943 1529 8977 1563
rect 8943 1461 8977 1495
rect 8943 1393 8977 1427
rect 8943 1325 8977 1359
rect 8943 1257 8977 1291
rect 8943 1189 8977 1223
rect 8943 1121 8977 1155
rect 8943 1053 8977 1087
rect 8943 985 8977 1019
rect 8943 917 8977 951
rect 8943 849 8977 883
rect 8943 781 8977 815
rect 8943 713 8977 747
rect 8943 645 8977 679
rect 8943 577 8977 611
rect 8943 509 8977 543
rect 8943 441 8977 475
rect 8943 373 8977 407
rect 8943 305 8977 339
rect 8943 237 8977 271
rect 8943 169 8977 203
rect 8943 101 8977 135
rect -317 -35 -283 -1
rect -92 -32 -58 2
rect 4093 -7 4127 27
rect 8943 33 8977 67
rect 8943 -35 8977 -1
rect -317 -103 -283 -69
rect -317 -171 -283 -137
rect -317 -239 -283 -205
rect -317 -307 -283 -273
rect -317 -375 -283 -341
rect -317 -443 -283 -409
rect -317 -511 -283 -477
rect -317 -579 -283 -545
rect -317 -647 -283 -613
rect -317 -715 -283 -681
rect -317 -783 -283 -749
rect -317 -851 -283 -817
rect -317 -919 -283 -885
rect -317 -987 -283 -953
rect -317 -1055 -283 -1021
rect -317 -1123 -283 -1089
rect -317 -1191 -283 -1157
rect -317 -1259 -283 -1225
rect -317 -1327 -283 -1293
rect -317 -1395 -283 -1361
rect -317 -1463 -283 -1429
rect -317 -1531 -283 -1497
rect -317 -1599 -283 -1565
rect -317 -1667 -283 -1633
rect -317 -1735 -283 -1701
rect -317 -1803 -283 -1769
rect -317 -1871 -283 -1837
rect -317 -1939 -283 -1905
rect -317 -2007 -283 -1973
rect -317 -2075 -283 -2041
rect -317 -2143 -283 -2109
rect -317 -2211 -283 -2177
rect -317 -2279 -283 -2245
rect -317 -2347 -283 -2313
rect -317 -2415 -283 -2381
rect -317 -2483 -283 -2449
rect -317 -2551 -283 -2517
rect -317 -2619 -283 -2585
rect -317 -2687 -283 -2653
rect -317 -2755 -283 -2721
rect -317 -2823 -283 -2789
rect -317 -2891 -283 -2857
rect -317 -2959 -283 -2925
rect -317 -3027 -283 -2993
rect -317 -3095 -283 -3061
rect -317 -3163 -283 -3129
rect -317 -3231 -283 -3197
rect -317 -3299 -283 -3265
rect -317 -3367 -283 -3333
rect -317 -3435 -283 -3401
rect -317 -3503 -283 -3469
rect -317 -3571 -283 -3537
rect -317 -3639 -283 -3605
rect -317 -3707 -283 -3673
rect -317 -3775 -283 -3741
rect -317 -3843 -283 -3809
rect -317 -3911 -283 -3877
rect -317 -3979 -283 -3945
rect -317 -4047 -283 -4013
rect -317 -4115 -283 -4081
rect -317 -4183 -283 -4149
rect -317 -4251 -283 -4217
rect -317 -4319 -283 -4285
rect -317 -4387 -283 -4353
rect -317 -4455 -283 -4421
rect -317 -4523 -283 -4489
rect -317 -4591 -283 -4557
rect -317 -4659 -283 -4625
rect -317 -4727 -283 -4693
rect -317 -4795 -283 -4761
rect -317 -4863 -283 -4829
rect -317 -4931 -283 -4897
rect -317 -4999 -283 -4965
rect -317 -5067 -283 -5033
rect -317 -5135 -283 -5101
rect 8943 -103 8977 -69
rect 8943 -171 8977 -137
rect 8943 -239 8977 -205
rect 8943 -307 8977 -273
rect 8943 -375 8977 -341
rect 8943 -443 8977 -409
rect 8943 -511 8977 -477
rect 8943 -579 8977 -545
rect 8943 -647 8977 -613
rect 8943 -715 8977 -681
rect 8943 -783 8977 -749
rect 8943 -851 8977 -817
rect 8943 -919 8977 -885
rect 8943 -987 8977 -953
rect 8943 -1055 8977 -1021
rect 8943 -1123 8977 -1089
rect 8943 -1191 8977 -1157
rect 8943 -1259 8977 -1225
rect 8943 -1327 8977 -1293
rect 8943 -1395 8977 -1361
rect 8943 -1463 8977 -1429
rect 8943 -1531 8977 -1497
rect 8943 -1599 8977 -1565
rect 8943 -1667 8977 -1633
rect 8943 -1735 8977 -1701
rect 8943 -1803 8977 -1769
rect 8943 -1871 8977 -1837
rect 8943 -1939 8977 -1905
rect 8943 -2007 8977 -1973
rect 8943 -2075 8977 -2041
rect 8943 -2143 8977 -2109
rect 8943 -2211 8977 -2177
rect 8943 -2279 8977 -2245
rect 8943 -2347 8977 -2313
rect 8943 -2415 8977 -2381
rect 8943 -2483 8977 -2449
rect 8943 -2551 8977 -2517
rect 8943 -2619 8977 -2585
rect 8943 -2687 8977 -2653
rect 8943 -2755 8977 -2721
rect 8943 -2823 8977 -2789
rect 8943 -2891 8977 -2857
rect 8943 -2959 8977 -2925
rect 8943 -3027 8977 -2993
rect 8943 -3095 8977 -3061
rect 8943 -3163 8977 -3129
rect 8943 -3231 8977 -3197
rect 8943 -3299 8977 -3265
rect 8943 -3367 8977 -3333
rect 8943 -3435 8977 -3401
rect 8943 -3503 8977 -3469
rect 8943 -3571 8977 -3537
rect 8943 -3639 8977 -3605
rect 8943 -3707 8977 -3673
rect 8943 -3775 8977 -3741
rect 8943 -3843 8977 -3809
rect 8943 -3911 8977 -3877
rect 8943 -3979 8977 -3945
rect 8943 -4047 8977 -4013
rect 8943 -4115 8977 -4081
rect 8943 -4183 8977 -4149
rect 8943 -4251 8977 -4217
rect 8943 -4319 8977 -4285
rect 8943 -4387 8977 -4353
rect 8943 -4455 8977 -4421
rect 8943 -4523 8977 -4489
rect 8943 -4591 8977 -4557
rect 8943 -4659 8977 -4625
rect 8943 -4727 8977 -4693
rect 8943 -4795 8977 -4761
rect 8943 -4863 8977 -4829
rect 8943 -4931 8977 -4897
rect 8943 -4999 8977 -4965
rect 8943 -5067 8977 -5033
rect 8943 -5135 8977 -5101
rect -243 -5217 -209 -5183
rect -175 -5217 -141 -5183
rect -107 -5217 -73 -5183
rect -39 -5217 -5 -5183
rect 29 -5217 63 -5183
rect 97 -5217 131 -5183
rect 165 -5217 199 -5183
rect 233 -5217 267 -5183
rect 301 -5217 335 -5183
rect 369 -5217 403 -5183
rect 437 -5217 471 -5183
rect 505 -5217 539 -5183
rect 573 -5217 607 -5183
rect 641 -5217 675 -5183
rect 709 -5217 743 -5183
rect 777 -5217 811 -5183
rect 845 -5217 879 -5183
rect 913 -5217 947 -5183
rect 981 -5217 1015 -5183
rect 1049 -5217 1083 -5183
rect 1117 -5217 1151 -5183
rect 1185 -5217 1219 -5183
rect 1253 -5217 1287 -5183
rect 1321 -5217 1355 -5183
rect 1389 -5217 1423 -5183
rect 1457 -5217 1491 -5183
rect 1525 -5217 1559 -5183
rect 1593 -5217 1627 -5183
rect 1661 -5217 1695 -5183
rect 1729 -5217 1763 -5183
rect 1797 -5217 1831 -5183
rect 1865 -5217 1899 -5183
rect 1933 -5217 1967 -5183
rect 2001 -5217 2035 -5183
rect 2069 -5217 2103 -5183
rect 2137 -5217 2171 -5183
rect 2205 -5217 2239 -5183
rect 2273 -5217 2307 -5183
rect 2341 -5217 2375 -5183
rect 2409 -5217 2443 -5183
rect 2477 -5217 2511 -5183
rect 2545 -5217 2579 -5183
rect 2613 -5217 2647 -5183
rect 2681 -5217 2715 -5183
rect 2749 -5217 2783 -5183
rect 2817 -5217 2851 -5183
rect 2885 -5217 2919 -5183
rect 2953 -5217 2987 -5183
rect 3021 -5217 3055 -5183
rect 3089 -5217 3123 -5183
rect 3157 -5217 3191 -5183
rect 3225 -5217 3259 -5183
rect 3293 -5217 3327 -5183
rect 3361 -5217 3395 -5183
rect 3429 -5217 3463 -5183
rect 3497 -5217 3531 -5183
rect 3565 -5217 3599 -5183
rect 3633 -5217 3667 -5183
rect 3701 -5217 3735 -5183
rect 3769 -5217 3803 -5183
rect 3837 -5217 3871 -5183
rect 3905 -5217 3939 -5183
rect 3973 -5217 4007 -5183
rect 4041 -5217 4075 -5183
rect 4109 -5217 4143 -5183
rect 4177 -5217 4211 -5183
rect 4245 -5217 4279 -5183
rect 4313 -5217 4347 -5183
rect 4381 -5217 4415 -5183
rect 4449 -5217 4483 -5183
rect 4517 -5217 4551 -5183
rect 4585 -5217 4619 -5183
rect 4653 -5217 4687 -5183
rect 4721 -5217 4755 -5183
rect 4789 -5217 4823 -5183
rect 4857 -5217 4891 -5183
rect 4925 -5217 4959 -5183
rect 4993 -5217 5027 -5183
rect 5061 -5217 5095 -5183
rect 5129 -5217 5163 -5183
rect 5197 -5217 5231 -5183
rect 5265 -5217 5299 -5183
rect 5333 -5217 5367 -5183
rect 5401 -5217 5435 -5183
rect 5469 -5217 5503 -5183
rect 5537 -5217 5571 -5183
rect 5605 -5217 5639 -5183
rect 5673 -5217 5707 -5183
rect 5741 -5217 5775 -5183
rect 5809 -5217 5843 -5183
rect 5877 -5217 5911 -5183
rect 5945 -5217 5979 -5183
rect 6013 -5217 6047 -5183
rect 6081 -5217 6115 -5183
rect 6149 -5217 6183 -5183
rect 6217 -5217 6251 -5183
rect 6285 -5217 6319 -5183
rect 6353 -5217 6387 -5183
rect 6421 -5217 6455 -5183
rect 6489 -5217 6523 -5183
rect 6557 -5217 6591 -5183
rect 6625 -5217 6659 -5183
rect 6693 -5217 6727 -5183
rect 6761 -5217 6795 -5183
rect 6829 -5217 6863 -5183
rect 6897 -5217 6931 -5183
rect 6965 -5217 6999 -5183
rect 7033 -5217 7067 -5183
rect 7101 -5217 7135 -5183
rect 7169 -5217 7203 -5183
rect 7237 -5217 7271 -5183
rect 7305 -5217 7339 -5183
rect 7373 -5217 7407 -5183
rect 7441 -5217 7475 -5183
rect 7509 -5217 7543 -5183
rect 7577 -5217 7611 -5183
rect 7645 -5217 7679 -5183
rect 7713 -5217 7747 -5183
rect 7781 -5217 7815 -5183
rect 7849 -5217 7883 -5183
rect 7917 -5217 7951 -5183
rect 7985 -5217 8019 -5183
rect 8053 -5217 8087 -5183
rect 8121 -5217 8155 -5183
rect 8189 -5217 8223 -5183
rect 8257 -5217 8291 -5183
rect 8325 -5217 8359 -5183
rect 8393 -5217 8427 -5183
rect 8461 -5217 8495 -5183
rect 8529 -5217 8563 -5183
rect 8597 -5217 8631 -5183
rect 8665 -5217 8699 -5183
rect 8733 -5217 8767 -5183
rect 8801 -5217 8835 -5183
rect 8869 -5217 8903 -5183
<< locali >>
rect -317 5283 -243 5317
rect -209 5283 -175 5317
rect -141 5283 -107 5317
rect -73 5283 -39 5317
rect -5 5283 29 5317
rect 63 5283 97 5317
rect 131 5283 165 5317
rect 199 5283 233 5317
rect 267 5283 301 5317
rect 335 5283 369 5317
rect 403 5283 437 5317
rect 471 5283 505 5317
rect 539 5283 573 5317
rect 607 5283 641 5317
rect 675 5283 709 5317
rect 743 5283 777 5317
rect 811 5283 845 5317
rect 879 5283 913 5317
rect 947 5283 981 5317
rect 1015 5283 1049 5317
rect 1083 5283 1117 5317
rect 1151 5283 1185 5317
rect 1219 5283 1253 5317
rect 1287 5283 1321 5317
rect 1355 5283 1389 5317
rect 1423 5283 1457 5317
rect 1491 5283 1525 5317
rect 1559 5283 1593 5317
rect 1627 5283 1661 5317
rect 1695 5283 1729 5317
rect 1763 5283 1797 5317
rect 1831 5283 1865 5317
rect 1899 5283 1933 5317
rect 1967 5283 2001 5317
rect 2035 5283 2069 5317
rect 2103 5283 2137 5317
rect 2171 5283 2205 5317
rect 2239 5283 2273 5317
rect 2307 5283 2341 5317
rect 2375 5283 2409 5317
rect 2443 5283 2477 5317
rect 2511 5283 2545 5317
rect 2579 5283 2613 5317
rect 2647 5283 2681 5317
rect 2715 5283 2749 5317
rect 2783 5283 2817 5317
rect 2851 5283 2885 5317
rect 2919 5283 2953 5317
rect 2987 5283 3021 5317
rect 3055 5283 3089 5317
rect 3123 5283 3157 5317
rect 3191 5283 3225 5317
rect 3259 5283 3293 5317
rect 3327 5283 3361 5317
rect 3395 5283 3429 5317
rect 3463 5283 3497 5317
rect 3531 5283 3565 5317
rect 3599 5283 3633 5317
rect 3667 5283 3701 5317
rect 3735 5283 3769 5317
rect 3803 5283 3837 5317
rect 3871 5283 3905 5317
rect 3939 5283 3973 5317
rect 4007 5283 4041 5317
rect 4075 5283 4109 5317
rect 4143 5283 4177 5317
rect 4211 5283 4245 5317
rect 4279 5283 4313 5317
rect 4347 5283 4381 5317
rect 4415 5283 4449 5317
rect 4483 5283 4517 5317
rect 4551 5283 4585 5317
rect 4619 5283 4653 5317
rect 4687 5283 4721 5317
rect 4755 5283 4789 5317
rect 4823 5283 4857 5317
rect 4891 5283 4925 5317
rect 4959 5283 4993 5317
rect 5027 5283 5061 5317
rect 5095 5283 5129 5317
rect 5163 5283 5197 5317
rect 5231 5283 5265 5317
rect 5299 5283 5333 5317
rect 5367 5283 5401 5317
rect 5435 5283 5469 5317
rect 5503 5283 5537 5317
rect 5571 5283 5605 5317
rect 5639 5283 5673 5317
rect 5707 5283 5741 5317
rect 5775 5283 5809 5317
rect 5843 5283 5877 5317
rect 5911 5283 5945 5317
rect 5979 5283 6013 5317
rect 6047 5283 6081 5317
rect 6115 5283 6149 5317
rect 6183 5283 6217 5317
rect 6251 5283 6285 5317
rect 6319 5283 6353 5317
rect 6387 5283 6421 5317
rect 6455 5283 6489 5317
rect 6523 5283 6557 5317
rect 6591 5283 6625 5317
rect 6659 5283 6693 5317
rect 6727 5283 6761 5317
rect 6795 5283 6829 5317
rect 6863 5283 6897 5317
rect 6931 5283 6965 5317
rect 6999 5283 7033 5317
rect 7067 5283 7101 5317
rect 7135 5283 7169 5317
rect 7203 5283 7237 5317
rect 7271 5283 7305 5317
rect 7339 5283 7373 5317
rect 7407 5283 7441 5317
rect 7475 5283 7509 5317
rect 7543 5283 7577 5317
rect 7611 5283 7645 5317
rect 7679 5283 7713 5317
rect 7747 5283 7781 5317
rect 7815 5283 7849 5317
rect 7883 5283 7917 5317
rect 7951 5283 7985 5317
rect 8019 5283 8053 5317
rect 8087 5283 8121 5317
rect 8155 5283 8189 5317
rect 8223 5283 8257 5317
rect 8291 5283 8325 5317
rect 8359 5283 8393 5317
rect 8427 5283 8461 5317
rect 8495 5283 8529 5317
rect 8563 5283 8597 5317
rect 8631 5283 8665 5317
rect 8699 5283 8733 5317
rect 8767 5283 8801 5317
rect 8835 5283 8869 5317
rect 8903 5283 8977 5317
rect -317 5235 -283 5283
rect -317 5167 -283 5201
rect -317 5099 -283 5133
rect -317 5031 -283 5065
rect -317 4963 -283 4997
rect -317 4895 -283 4929
rect -317 4827 -283 4861
rect -317 4759 -283 4793
rect -317 4691 -283 4725
rect -317 4623 -283 4657
rect -317 4555 -283 4589
rect -317 4487 -283 4521
rect -317 4419 -283 4453
rect -317 4351 -283 4385
rect -317 4283 -283 4317
rect -317 4215 -283 4249
rect -317 4147 -283 4181
rect -317 4079 -283 4113
rect -317 4011 -283 4045
rect -317 3943 -283 3977
rect -317 3875 -283 3909
rect -317 3807 -283 3841
rect -317 3739 -283 3773
rect -317 3671 -283 3705
rect -317 3603 -283 3637
rect -317 3535 -283 3569
rect -317 3467 -283 3501
rect -317 3399 -283 3433
rect -317 3331 -283 3365
rect -317 3263 -283 3297
rect -317 3195 -283 3229
rect -317 3127 -283 3161
rect -317 3059 -283 3093
rect -317 2991 -283 3025
rect -317 2923 -283 2957
rect -317 2855 -283 2889
rect -317 2787 -283 2821
rect -317 2719 -283 2753
rect -317 2651 -283 2685
rect -317 2583 -283 2617
rect -317 2515 -283 2549
rect -317 2447 -283 2481
rect -317 2379 -283 2413
rect -317 2311 -283 2345
rect -317 2243 -283 2277
rect -317 2175 -283 2209
rect -317 2107 -283 2141
rect -317 2039 -283 2073
rect -317 1971 -283 2005
rect -317 1903 -283 1937
rect -317 1835 -283 1869
rect -317 1767 -283 1801
rect -317 1699 -283 1733
rect -317 1631 -283 1665
rect -317 1563 -283 1597
rect -317 1495 -283 1529
rect -317 1427 -283 1461
rect -317 1359 -283 1393
rect -317 1291 -283 1325
rect -317 1223 -283 1257
rect -317 1155 -283 1189
rect -317 1087 -283 1121
rect -317 1019 -283 1053
rect -317 951 -283 985
rect -317 883 -283 917
rect -317 815 -283 849
rect -317 747 -283 781
rect -317 679 -283 713
rect -317 611 -283 645
rect -317 543 -283 577
rect -317 475 -283 509
rect -317 407 -283 441
rect -317 339 -283 373
rect -317 271 -283 305
rect -317 203 -283 237
rect -317 135 -283 169
rect -317 67 -283 101
rect 8943 5235 8977 5283
rect 8943 5167 8977 5201
rect 8943 5099 8977 5133
rect 8943 5031 8977 5065
rect 8943 4963 8977 4997
rect 8943 4895 8977 4929
rect 8943 4827 8977 4861
rect 8943 4759 8977 4793
rect 8943 4691 8977 4725
rect 8943 4623 8977 4657
rect 8943 4555 8977 4589
rect 8943 4487 8977 4521
rect 8943 4419 8977 4453
rect 8943 4351 8977 4385
rect 8943 4283 8977 4317
rect 8943 4215 8977 4249
rect 8943 4147 8977 4181
rect 8943 4079 8977 4113
rect 8943 4011 8977 4045
rect 8943 3943 8977 3977
rect 8943 3875 8977 3909
rect 8943 3807 8977 3841
rect 8943 3739 8977 3773
rect 8943 3671 8977 3705
rect 8943 3603 8977 3637
rect 8943 3535 8977 3569
rect 8943 3467 8977 3501
rect 8943 3399 8977 3433
rect 8943 3331 8977 3365
rect 8943 3263 8977 3297
rect 8943 3195 8977 3229
rect 8943 3127 8977 3161
rect 8943 3059 8977 3093
rect 8943 2991 8977 3025
rect 8943 2923 8977 2957
rect 8943 2855 8977 2889
rect 8943 2787 8977 2821
rect 8943 2719 8977 2753
rect 8943 2651 8977 2685
rect 8943 2583 8977 2617
rect 8943 2515 8977 2549
rect 8943 2447 8977 2481
rect 8943 2379 8977 2413
rect 8943 2311 8977 2345
rect 8943 2243 8977 2277
rect 8943 2175 8977 2209
rect 8943 2107 8977 2141
rect 8943 2039 8977 2073
rect 8943 1971 8977 2005
rect 8943 1903 8977 1937
rect 8943 1835 8977 1869
rect 8943 1767 8977 1801
rect 8943 1699 8977 1733
rect 8943 1631 8977 1665
rect 8943 1563 8977 1597
rect 8943 1495 8977 1529
rect 8943 1427 8977 1461
rect 8943 1359 8977 1393
rect 8943 1291 8977 1325
rect 8943 1223 8977 1257
rect 8943 1155 8977 1189
rect 8943 1087 8977 1121
rect 8943 1019 8977 1053
rect 8943 951 8977 985
rect 8943 883 8977 917
rect 8943 815 8977 849
rect 8943 747 8977 781
rect 8943 679 8977 713
rect 8943 611 8977 645
rect 8943 543 8977 577
rect 8943 475 8977 509
rect 8943 407 8977 441
rect 8943 339 8977 373
rect 8943 271 8977 305
rect 8943 203 8977 237
rect 8943 135 8977 169
rect 8943 67 8977 101
rect -317 -1 -283 33
rect 4090 27 4130 46
rect -317 -69 -283 -35
rect -100 2 -50 26
rect -100 -32 -92 2
rect -58 -32 -50 2
rect 4090 -7 4093 27
rect 4127 -7 4130 27
rect 4090 -26 4130 -7
rect 8943 -1 8977 33
rect -100 -56 -50 -32
rect -317 -137 -283 -103
rect -317 -205 -283 -171
rect -317 -273 -283 -239
rect -317 -341 -283 -307
rect -317 -409 -283 -375
rect -317 -477 -283 -443
rect -317 -545 -283 -511
rect -317 -613 -283 -579
rect -317 -681 -283 -647
rect -317 -749 -283 -715
rect -317 -817 -283 -783
rect -317 -885 -283 -851
rect -317 -953 -283 -919
rect -317 -1021 -283 -987
rect -317 -1089 -283 -1055
rect -317 -1157 -283 -1123
rect -317 -1225 -283 -1191
rect -317 -1293 -283 -1259
rect -317 -1361 -283 -1327
rect -317 -1429 -283 -1395
rect -317 -1497 -283 -1463
rect -317 -1565 -283 -1531
rect -317 -1633 -283 -1599
rect -317 -1701 -283 -1667
rect -317 -1769 -283 -1735
rect -317 -1837 -283 -1803
rect -317 -1905 -283 -1871
rect -317 -1973 -283 -1939
rect -317 -2041 -283 -2007
rect -317 -2109 -283 -2075
rect -317 -2177 -283 -2143
rect -317 -2245 -283 -2211
rect -317 -2313 -283 -2279
rect -317 -2381 -283 -2347
rect -317 -2449 -283 -2415
rect -317 -2517 -283 -2483
rect -317 -2585 -283 -2551
rect -317 -2653 -283 -2619
rect -317 -2721 -283 -2687
rect -317 -2789 -283 -2755
rect -317 -2857 -283 -2823
rect -317 -2925 -283 -2891
rect -317 -2993 -283 -2959
rect -317 -3061 -283 -3027
rect -317 -3129 -283 -3095
rect -317 -3197 -283 -3163
rect -317 -3265 -283 -3231
rect -317 -3333 -283 -3299
rect -317 -3401 -283 -3367
rect -317 -3469 -283 -3435
rect -317 -3537 -283 -3503
rect -317 -3605 -283 -3571
rect -317 -3673 -283 -3639
rect -317 -3741 -283 -3707
rect -317 -3809 -283 -3775
rect -317 -3877 -283 -3843
rect -317 -3945 -283 -3911
rect -317 -4013 -283 -3979
rect -317 -4081 -283 -4047
rect -317 -4149 -283 -4115
rect -317 -4217 -283 -4183
rect -317 -4285 -283 -4251
rect -317 -4353 -283 -4319
rect -317 -4421 -283 -4387
rect -317 -4489 -283 -4455
rect -317 -4557 -283 -4523
rect -317 -4625 -283 -4591
rect -317 -4693 -283 -4659
rect -317 -4761 -283 -4727
rect -317 -4829 -283 -4795
rect -317 -4897 -283 -4863
rect -317 -4965 -283 -4931
rect -317 -5033 -283 -4999
rect -317 -5101 -283 -5067
rect -317 -5183 -283 -5135
rect 8943 -69 8977 -35
rect 8943 -137 8977 -103
rect 8943 -205 8977 -171
rect 8943 -273 8977 -239
rect 8943 -341 8977 -307
rect 8943 -409 8977 -375
rect 8943 -477 8977 -443
rect 8943 -545 8977 -511
rect 8943 -613 8977 -579
rect 8943 -681 8977 -647
rect 8943 -749 8977 -715
rect 8943 -817 8977 -783
rect 8943 -885 8977 -851
rect 8943 -953 8977 -919
rect 8943 -1021 8977 -987
rect 8943 -1089 8977 -1055
rect 8943 -1157 8977 -1123
rect 8943 -1225 8977 -1191
rect 8943 -1293 8977 -1259
rect 8943 -1361 8977 -1327
rect 8943 -1429 8977 -1395
rect 8943 -1497 8977 -1463
rect 8943 -1565 8977 -1531
rect 8943 -1633 8977 -1599
rect 8943 -1701 8977 -1667
rect 8943 -1769 8977 -1735
rect 8943 -1837 8977 -1803
rect 8943 -1905 8977 -1871
rect 8943 -1973 8977 -1939
rect 8943 -2041 8977 -2007
rect 8943 -2109 8977 -2075
rect 8943 -2177 8977 -2143
rect 8943 -2245 8977 -2211
rect 8943 -2313 8977 -2279
rect 8943 -2381 8977 -2347
rect 8943 -2449 8977 -2415
rect 8943 -2517 8977 -2483
rect 8943 -2585 8977 -2551
rect 8943 -2653 8977 -2619
rect 8943 -2721 8977 -2687
rect 8943 -2789 8977 -2755
rect 8943 -2857 8977 -2823
rect 8943 -2925 8977 -2891
rect 8943 -2993 8977 -2959
rect 8943 -3061 8977 -3027
rect 8943 -3129 8977 -3095
rect 8943 -3197 8977 -3163
rect 8943 -3265 8977 -3231
rect 8943 -3333 8977 -3299
rect 8943 -3401 8977 -3367
rect 8943 -3469 8977 -3435
rect 8943 -3537 8977 -3503
rect 8943 -3605 8977 -3571
rect 8943 -3673 8977 -3639
rect 8943 -3741 8977 -3707
rect 8943 -3809 8977 -3775
rect 8943 -3877 8977 -3843
rect 8943 -3945 8977 -3911
rect 8943 -4013 8977 -3979
rect 8943 -4081 8977 -4047
rect 8943 -4149 8977 -4115
rect 8943 -4217 8977 -4183
rect 8943 -4285 8977 -4251
rect 8943 -4353 8977 -4319
rect 8943 -4421 8977 -4387
rect 8943 -4489 8977 -4455
rect 8943 -4557 8977 -4523
rect 8943 -4625 8977 -4591
rect 8943 -4693 8977 -4659
rect 8943 -4761 8977 -4727
rect 8943 -4829 8977 -4795
rect 8943 -4897 8977 -4863
rect 8943 -4965 8977 -4931
rect 8943 -5033 8977 -4999
rect 8943 -5101 8977 -5067
rect 8943 -5183 8977 -5135
rect -317 -5217 -243 -5183
rect -209 -5217 -175 -5183
rect -141 -5217 -107 -5183
rect -73 -5217 -39 -5183
rect -5 -5217 29 -5183
rect 63 -5217 97 -5183
rect 131 -5217 165 -5183
rect 199 -5217 233 -5183
rect 267 -5217 301 -5183
rect 335 -5217 369 -5183
rect 403 -5217 437 -5183
rect 471 -5217 505 -5183
rect 539 -5217 573 -5183
rect 607 -5217 641 -5183
rect 675 -5217 709 -5183
rect 743 -5217 777 -5183
rect 811 -5217 845 -5183
rect 879 -5217 913 -5183
rect 947 -5217 981 -5183
rect 1015 -5217 1049 -5183
rect 1083 -5217 1117 -5183
rect 1151 -5217 1185 -5183
rect 1219 -5217 1253 -5183
rect 1287 -5217 1321 -5183
rect 1355 -5217 1389 -5183
rect 1423 -5217 1457 -5183
rect 1491 -5217 1525 -5183
rect 1559 -5217 1593 -5183
rect 1627 -5217 1661 -5183
rect 1695 -5217 1729 -5183
rect 1763 -5217 1797 -5183
rect 1831 -5217 1865 -5183
rect 1899 -5217 1933 -5183
rect 1967 -5217 2001 -5183
rect 2035 -5217 2069 -5183
rect 2103 -5217 2137 -5183
rect 2171 -5217 2205 -5183
rect 2239 -5217 2273 -5183
rect 2307 -5217 2341 -5183
rect 2375 -5217 2409 -5183
rect 2443 -5217 2477 -5183
rect 2511 -5217 2545 -5183
rect 2579 -5217 2613 -5183
rect 2647 -5217 2681 -5183
rect 2715 -5217 2749 -5183
rect 2783 -5217 2817 -5183
rect 2851 -5217 2885 -5183
rect 2919 -5217 2953 -5183
rect 2987 -5217 3021 -5183
rect 3055 -5217 3089 -5183
rect 3123 -5217 3157 -5183
rect 3191 -5217 3225 -5183
rect 3259 -5217 3293 -5183
rect 3327 -5217 3361 -5183
rect 3395 -5217 3429 -5183
rect 3463 -5217 3497 -5183
rect 3531 -5217 3565 -5183
rect 3599 -5217 3633 -5183
rect 3667 -5217 3701 -5183
rect 3735 -5217 3769 -5183
rect 3803 -5217 3837 -5183
rect 3871 -5217 3905 -5183
rect 3939 -5217 3973 -5183
rect 4007 -5217 4041 -5183
rect 4075 -5217 4109 -5183
rect 4143 -5217 4177 -5183
rect 4211 -5217 4245 -5183
rect 4279 -5217 4313 -5183
rect 4347 -5217 4381 -5183
rect 4415 -5217 4449 -5183
rect 4483 -5217 4517 -5183
rect 4551 -5217 4585 -5183
rect 4619 -5217 4653 -5183
rect 4687 -5217 4721 -5183
rect 4755 -5217 4789 -5183
rect 4823 -5217 4857 -5183
rect 4891 -5217 4925 -5183
rect 4959 -5217 4993 -5183
rect 5027 -5217 5061 -5183
rect 5095 -5217 5129 -5183
rect 5163 -5217 5197 -5183
rect 5231 -5217 5265 -5183
rect 5299 -5217 5333 -5183
rect 5367 -5217 5401 -5183
rect 5435 -5217 5469 -5183
rect 5503 -5217 5537 -5183
rect 5571 -5217 5605 -5183
rect 5639 -5217 5673 -5183
rect 5707 -5217 5741 -5183
rect 5775 -5217 5809 -5183
rect 5843 -5217 5877 -5183
rect 5911 -5217 5945 -5183
rect 5979 -5217 6013 -5183
rect 6047 -5217 6081 -5183
rect 6115 -5217 6149 -5183
rect 6183 -5217 6217 -5183
rect 6251 -5217 6285 -5183
rect 6319 -5217 6353 -5183
rect 6387 -5217 6421 -5183
rect 6455 -5217 6489 -5183
rect 6523 -5217 6557 -5183
rect 6591 -5217 6625 -5183
rect 6659 -5217 6693 -5183
rect 6727 -5217 6761 -5183
rect 6795 -5217 6829 -5183
rect 6863 -5217 6897 -5183
rect 6931 -5217 6965 -5183
rect 6999 -5217 7033 -5183
rect 7067 -5217 7101 -5183
rect 7135 -5217 7169 -5183
rect 7203 -5217 7237 -5183
rect 7271 -5217 7305 -5183
rect 7339 -5217 7373 -5183
rect 7407 -5217 7441 -5183
rect 7475 -5217 7509 -5183
rect 7543 -5217 7577 -5183
rect 7611 -5217 7645 -5183
rect 7679 -5217 7713 -5183
rect 7747 -5217 7781 -5183
rect 7815 -5217 7849 -5183
rect 7883 -5217 7917 -5183
rect 7951 -5217 7985 -5183
rect 8019 -5217 8053 -5183
rect 8087 -5217 8121 -5183
rect 8155 -5217 8189 -5183
rect 8223 -5217 8257 -5183
rect 8291 -5217 8325 -5183
rect 8359 -5217 8393 -5183
rect 8427 -5217 8461 -5183
rect 8495 -5217 8529 -5183
rect 8563 -5217 8597 -5183
rect 8631 -5217 8665 -5183
rect 8699 -5217 8733 -5183
rect 8767 -5217 8801 -5183
rect 8835 -5217 8869 -5183
rect 8903 -5217 8977 -5183
<< viali >>
rect -92 -32 -58 2
rect 4093 -7 4127 27
<< metal1 >>
rect 10 5010 220 5510
rect 1500 5160 1640 5510
rect 8750 5086 8910 5100
rect 8750 5034 8764 5086
rect 8816 5034 8844 5086
rect 8896 5034 8910 5086
rect 8750 5020 8910 5034
rect 10 4900 210 5010
rect 10 4690 220 4900
rect 2130 4766 2290 4770
rect 2130 4714 2144 4766
rect 2196 4714 2224 4766
rect 2276 4714 2290 4766
rect 2130 4710 2290 4714
rect 10 4680 2100 4690
rect 10 4630 2200 4680
rect 240 4430 2200 4630
rect 20 4426 2200 4430
rect 20 4374 1934 4426
rect 1986 4374 2014 4426
rect 2066 4374 2200 4426
rect 20 4370 2200 4374
rect 20 4250 300 4370
rect 420 4306 570 4310
rect 420 4254 437 4306
rect 489 4254 501 4306
rect 553 4254 570 4306
rect 420 4250 570 4254
rect 800 4306 950 4310
rect 800 4254 817 4306
rect 869 4254 881 4306
rect 933 4254 950 4306
rect 800 4250 950 4254
rect 1180 4306 1330 4310
rect 1180 4254 1197 4306
rect 1249 4254 1261 4306
rect 1313 4254 1330 4306
rect 1180 4250 1330 4254
rect 1560 4306 1710 4310
rect 1560 4254 1577 4306
rect 1629 4254 1641 4306
rect 1693 4254 1710 4306
rect 1560 4250 1710 4254
rect 1940 4306 2090 4310
rect 1940 4254 1957 4306
rect 2009 4254 2021 4306
rect 2073 4254 2090 4306
rect 1940 4250 2090 4254
rect -110 2326 -30 2330
rect -110 2274 -96 2326
rect -44 2274 -30 2326
rect -110 2246 -30 2274
rect 240 2250 300 4250
rect 600 3526 680 3540
rect 600 3474 614 3526
rect 666 3474 680 3526
rect 600 3436 680 3474
rect 600 3384 614 3436
rect 666 3384 680 3436
rect 600 3346 680 3384
rect 600 3294 614 3346
rect 666 3294 680 3346
rect 600 3256 680 3294
rect 600 3204 614 3256
rect 666 3204 680 3256
rect 600 3166 680 3204
rect 600 3114 614 3166
rect 666 3114 680 3166
rect 600 3076 680 3114
rect 600 3024 614 3076
rect 666 3024 680 3076
rect 600 3010 680 3024
rect 980 3526 1060 3540
rect 980 3474 994 3526
rect 1046 3474 1060 3526
rect 980 3436 1060 3474
rect 980 3384 994 3436
rect 1046 3384 1060 3436
rect 980 3346 1060 3384
rect 980 3294 994 3346
rect 1046 3294 1060 3346
rect 980 3256 1060 3294
rect 980 3204 994 3256
rect 1046 3204 1060 3256
rect 980 3166 1060 3204
rect 980 3114 994 3166
rect 1046 3114 1060 3166
rect 980 3076 1060 3114
rect 980 3024 994 3076
rect 1046 3024 1060 3076
rect 980 3010 1060 3024
rect 1360 3526 1440 3540
rect 1360 3474 1374 3526
rect 1426 3474 1440 3526
rect 1360 3436 1440 3474
rect 1360 3384 1374 3436
rect 1426 3384 1440 3436
rect 1360 3346 1440 3384
rect 1360 3294 1374 3346
rect 1426 3294 1440 3346
rect 1360 3256 1440 3294
rect 1360 3204 1374 3256
rect 1426 3204 1440 3256
rect 1360 3166 1440 3204
rect 1360 3114 1374 3166
rect 1426 3114 1440 3166
rect 1360 3076 1440 3114
rect 1360 3024 1374 3076
rect 1426 3024 1440 3076
rect 1360 3010 1440 3024
rect 1740 3526 1820 3540
rect 1740 3474 1754 3526
rect 1806 3474 1820 3526
rect 1740 3436 1820 3474
rect 1740 3384 1754 3436
rect 1806 3384 1820 3436
rect 1740 3346 1820 3384
rect 1740 3294 1754 3346
rect 1806 3294 1820 3346
rect 1740 3256 1820 3294
rect 1740 3204 1754 3256
rect 1806 3204 1820 3256
rect 1740 3166 1820 3204
rect 1740 3114 1754 3166
rect 1806 3114 1820 3166
rect 1740 3076 1820 3114
rect 1740 3024 1754 3076
rect 1806 3024 1820 3076
rect 1740 3010 1820 3024
rect 2120 3526 2200 3540
rect 2120 3474 2134 3526
rect 2186 3474 2200 3526
rect 2120 3436 2200 3474
rect 2120 3384 2134 3436
rect 2186 3384 2200 3436
rect 2120 3346 2200 3384
rect 2120 3294 2134 3346
rect 2186 3294 2200 3346
rect 2120 3256 2200 3294
rect 2120 3204 2134 3256
rect 2186 3204 2200 3256
rect 2120 3166 2200 3204
rect 2120 3114 2134 3166
rect 2186 3114 2200 3166
rect 2120 3076 2200 3114
rect 2120 3024 2134 3076
rect 2186 3024 2200 3076
rect 2120 3010 2200 3024
rect 2230 2250 2290 4710
rect 2320 4426 8660 4690
rect 2320 4374 2334 4426
rect 2386 4374 2434 4426
rect 2486 4374 8660 4426
rect 2320 4370 8660 4374
rect 2320 4306 2470 4310
rect 2320 4254 2337 4306
rect 2389 4254 2401 4306
rect 2453 4254 2470 4306
rect 2320 4250 2470 4254
rect 2700 4306 2850 4310
rect 2700 4254 2717 4306
rect 2769 4254 2781 4306
rect 2833 4254 2850 4306
rect 2700 4250 2850 4254
rect 3080 4306 3230 4310
rect 3080 4254 3097 4306
rect 3149 4254 3161 4306
rect 3213 4254 3230 4306
rect 3080 4250 3230 4254
rect 3460 4306 3610 4310
rect 3460 4254 3477 4306
rect 3529 4254 3541 4306
rect 3593 4254 3610 4306
rect 3460 4250 3610 4254
rect 3840 4306 3990 4310
rect 3840 4254 3857 4306
rect 3909 4254 3921 4306
rect 3973 4254 3990 4306
rect 3840 4250 3990 4254
rect 4200 4250 4480 4370
rect 2500 3526 2580 3540
rect 2500 3474 2514 3526
rect 2566 3474 2580 3526
rect 2500 3436 2580 3474
rect 2500 3384 2514 3436
rect 2566 3384 2580 3436
rect 2500 3346 2580 3384
rect 2500 3294 2514 3346
rect 2566 3294 2580 3346
rect 2500 3256 2580 3294
rect 2500 3204 2514 3256
rect 2566 3204 2580 3256
rect 2500 3166 2580 3204
rect 2500 3114 2514 3166
rect 2566 3114 2580 3166
rect 2500 3076 2580 3114
rect 2500 3024 2514 3076
rect 2566 3024 2580 3076
rect 2500 3010 2580 3024
rect 2880 3526 2960 3540
rect 2880 3474 2894 3526
rect 2946 3474 2960 3526
rect 2880 3436 2960 3474
rect 2880 3384 2894 3436
rect 2946 3384 2960 3436
rect 2880 3346 2960 3384
rect 2880 3294 2894 3346
rect 2946 3294 2960 3346
rect 2880 3256 2960 3294
rect 2880 3204 2894 3256
rect 2946 3204 2960 3256
rect 2880 3166 2960 3204
rect 2880 3114 2894 3166
rect 2946 3114 2960 3166
rect 2880 3076 2960 3114
rect 2880 3024 2894 3076
rect 2946 3024 2960 3076
rect 2880 3010 2960 3024
rect 3260 3526 3340 3540
rect 3260 3474 3274 3526
rect 3326 3474 3340 3526
rect 3260 3436 3340 3474
rect 3260 3384 3274 3436
rect 3326 3384 3340 3436
rect 3260 3346 3340 3384
rect 3260 3294 3274 3346
rect 3326 3294 3340 3346
rect 3260 3256 3340 3294
rect 3260 3204 3274 3256
rect 3326 3204 3340 3256
rect 3260 3166 3340 3204
rect 3260 3114 3274 3166
rect 3326 3114 3340 3166
rect 3260 3076 3340 3114
rect 3260 3024 3274 3076
rect 3326 3024 3340 3076
rect 3260 3010 3340 3024
rect 3640 3526 3720 3540
rect 3640 3474 3654 3526
rect 3706 3474 3720 3526
rect 3640 3436 3720 3474
rect 3640 3384 3654 3436
rect 3706 3384 3720 3436
rect 3640 3346 3720 3384
rect 3640 3294 3654 3346
rect 3706 3294 3720 3346
rect 3640 3256 3720 3294
rect 3640 3204 3654 3256
rect 3706 3204 3720 3256
rect 3640 3166 3720 3204
rect 3640 3114 3654 3166
rect 3706 3114 3720 3166
rect 3640 3076 3720 3114
rect 3640 3024 3654 3076
rect 3706 3024 3720 3076
rect 3640 3010 3720 3024
rect 4020 3526 4100 3540
rect 4020 3474 4034 3526
rect 4086 3474 4100 3526
rect 4020 3436 4100 3474
rect 4020 3384 4034 3436
rect 4086 3384 4100 3436
rect 4020 3346 4100 3384
rect 4020 3294 4034 3346
rect 4086 3294 4100 3346
rect 4020 3256 4100 3294
rect 4020 3204 4034 3256
rect 4086 3204 4100 3256
rect 4020 3166 4100 3204
rect 4020 3114 4034 3166
rect 4086 3114 4100 3166
rect 4020 3076 4100 3114
rect 4020 3024 4034 3076
rect 4086 3024 4100 3076
rect 4020 3010 4100 3024
rect 4420 2250 4480 4250
rect -110 2194 -96 2246
rect -44 2194 -30 2246
rect -110 1796 -30 2194
rect 10 2070 300 2250
rect 420 2246 570 2250
rect 420 2194 437 2246
rect 489 2194 501 2246
rect 553 2194 570 2246
rect 420 2190 570 2194
rect 800 2246 950 2250
rect 800 2194 817 2246
rect 869 2194 881 2246
rect 933 2194 950 2246
rect 800 2190 950 2194
rect 1180 2246 1330 2250
rect 1180 2194 1197 2246
rect 1249 2194 1261 2246
rect 1313 2194 1330 2246
rect 1180 2190 1330 2194
rect 1560 2246 1710 2250
rect 1560 2194 1577 2246
rect 1629 2194 1641 2246
rect 1693 2194 1710 2246
rect 1560 2190 1710 2194
rect 1940 2246 2090 2250
rect 1940 2194 1957 2246
rect 2009 2194 2021 2246
rect 2073 2194 2090 2246
rect 1940 2190 2090 2194
rect 2230 2246 2470 2250
rect 2230 2194 2337 2246
rect 2389 2194 2401 2246
rect 2453 2194 2470 2246
rect 2230 2190 2470 2194
rect 2700 2246 2850 2250
rect 2700 2194 2717 2246
rect 2769 2194 2781 2246
rect 2833 2194 2850 2246
rect 2700 2190 2850 2194
rect 3080 2246 3230 2250
rect 3080 2194 3097 2246
rect 3149 2194 3161 2246
rect 3213 2194 3230 2246
rect 3080 2190 3230 2194
rect 3460 2246 3610 2250
rect 3460 2194 3477 2246
rect 3529 2194 3541 2246
rect 3593 2194 3610 2246
rect 3460 2190 3610 2194
rect 3840 2246 3990 2250
rect 3840 2194 3857 2246
rect 3909 2194 3921 2246
rect 3973 2194 3990 2246
rect 3840 2190 3990 2194
rect 4130 2190 4480 2250
rect 4510 4316 4700 4330
rect 4510 4264 4524 4316
rect 4576 4311 4700 4316
rect 4576 4264 4614 4311
rect 4510 4259 4614 4264
rect 4666 4310 4700 4311
rect 4666 4306 4750 4310
rect 4666 4259 4685 4306
rect 4510 4254 4685 4259
rect 4737 4254 4750 4306
rect 4510 4250 4750 4254
rect 4980 4306 5130 4310
rect 4980 4254 4997 4306
rect 5049 4254 5061 4306
rect 5113 4254 5130 4306
rect 4980 4250 5130 4254
rect 5360 4306 5510 4310
rect 5360 4254 5377 4306
rect 5429 4254 5441 4306
rect 5493 4254 5510 4306
rect 5360 4250 5510 4254
rect 5740 4306 5890 4310
rect 5740 4254 5757 4306
rect 5809 4254 5821 4306
rect 5873 4254 5890 4306
rect 5740 4250 5890 4254
rect 6120 4306 6270 4310
rect 6120 4254 6137 4306
rect 6189 4254 6201 4306
rect 6253 4254 6270 4306
rect 6120 4250 6270 4254
rect 6500 4306 6650 4310
rect 6500 4254 6517 4306
rect 6569 4254 6581 4306
rect 6633 4254 6650 4306
rect 6500 4250 6650 4254
rect 6880 4306 7030 4310
rect 6880 4254 6897 4306
rect 6949 4254 6961 4306
rect 7013 4254 7030 4306
rect 6880 4250 7030 4254
rect 7260 4306 7410 4310
rect 7260 4254 7277 4306
rect 7329 4254 7341 4306
rect 7393 4254 7410 4306
rect 7260 4250 7410 4254
rect 7640 4306 7790 4310
rect 7640 4254 7657 4306
rect 7709 4254 7721 4306
rect 7773 4254 7790 4306
rect 7640 4250 7790 4254
rect 8020 4306 8170 4310
rect 8020 4254 8037 4306
rect 8089 4254 8101 4306
rect 8153 4254 8170 4306
rect 8020 4250 8170 4254
rect 8370 4250 8660 4370
rect 420 2126 570 2130
rect 420 2074 437 2126
rect 489 2074 501 2126
rect 553 2074 570 2126
rect 420 2070 570 2074
rect 800 2126 950 2130
rect 800 2074 817 2126
rect 869 2074 881 2126
rect 933 2074 950 2126
rect 800 2070 950 2074
rect 1180 2126 1330 2130
rect 1180 2074 1197 2126
rect 1249 2074 1261 2126
rect 1313 2074 1330 2126
rect 1180 2070 1330 2074
rect 1560 2126 1710 2130
rect 1560 2074 1577 2126
rect 1629 2074 1641 2126
rect 1693 2074 1710 2126
rect 1560 2070 1710 2074
rect 1940 2126 2090 2130
rect 1940 2074 1957 2126
rect 2009 2074 2021 2126
rect 2073 2074 2090 2126
rect 1940 2070 2090 2074
rect -110 1744 -96 1796
rect -44 1744 -30 1796
rect -110 1706 -30 1744
rect -110 1654 -96 1706
rect -44 1654 -30 1706
rect -110 1640 -30 1654
rect 240 70 300 2070
rect 600 1376 680 1390
rect 600 1324 614 1376
rect 666 1324 680 1376
rect 600 1286 680 1324
rect 600 1234 614 1286
rect 666 1234 680 1286
rect 600 1196 680 1234
rect 600 1144 614 1196
rect 666 1144 680 1196
rect 600 1106 680 1144
rect 600 1054 614 1106
rect 666 1054 680 1106
rect 600 1016 680 1054
rect 600 964 614 1016
rect 666 964 680 1016
rect 600 926 680 964
rect 600 874 614 926
rect 666 874 680 926
rect 600 860 680 874
rect 980 1376 1060 1390
rect 980 1324 994 1376
rect 1046 1324 1060 1376
rect 980 1286 1060 1324
rect 980 1234 994 1286
rect 1046 1234 1060 1286
rect 980 1196 1060 1234
rect 980 1144 994 1196
rect 1046 1144 1060 1196
rect 980 1106 1060 1144
rect 980 1054 994 1106
rect 1046 1054 1060 1106
rect 980 1016 1060 1054
rect 980 964 994 1016
rect 1046 964 1060 1016
rect 980 926 1060 964
rect 980 874 994 926
rect 1046 874 1060 926
rect 980 860 1060 874
rect 1360 1376 1440 1390
rect 1360 1324 1374 1376
rect 1426 1324 1440 1376
rect 1360 1286 1440 1324
rect 1360 1234 1374 1286
rect 1426 1234 1440 1286
rect 1360 1196 1440 1234
rect 1360 1144 1374 1196
rect 1426 1144 1440 1196
rect 1360 1106 1440 1144
rect 1360 1054 1374 1106
rect 1426 1054 1440 1106
rect 1360 1016 1440 1054
rect 1360 964 1374 1016
rect 1426 964 1440 1016
rect 1360 926 1440 964
rect 1360 874 1374 926
rect 1426 874 1440 926
rect 1360 860 1440 874
rect 1740 1376 1820 1390
rect 1740 1324 1754 1376
rect 1806 1324 1820 1376
rect 1740 1286 1820 1324
rect 1740 1234 1754 1286
rect 1806 1234 1820 1286
rect 1740 1196 1820 1234
rect 1740 1144 1754 1196
rect 1806 1144 1820 1196
rect 1740 1106 1820 1144
rect 1740 1054 1754 1106
rect 1806 1054 1820 1106
rect 1740 1016 1820 1054
rect 1740 964 1754 1016
rect 1806 964 1820 1016
rect 1740 926 1820 964
rect 1740 874 1754 926
rect 1806 874 1820 926
rect 1740 860 1820 874
rect 2120 1376 2200 1390
rect 2120 1324 2134 1376
rect 2186 1324 2200 1376
rect 2120 1286 2200 1324
rect 2120 1234 2134 1286
rect 2186 1234 2200 1286
rect 2120 1196 2200 1234
rect 2120 1144 2134 1196
rect 2186 1144 2200 1196
rect 2120 1106 2200 1144
rect 2120 1054 2134 1106
rect 2186 1054 2200 1106
rect 2120 1016 2200 1054
rect 2120 964 2134 1016
rect 2186 964 2200 1016
rect 2120 926 2200 964
rect 2120 874 2134 926
rect 2186 874 2200 926
rect 2120 860 2200 874
rect 2230 70 2290 2190
rect 2320 2126 2470 2130
rect 2320 2074 2337 2126
rect 2389 2074 2401 2126
rect 2453 2074 2470 2126
rect 2320 2070 2470 2074
rect 2700 2126 2850 2130
rect 2700 2074 2717 2126
rect 2769 2074 2781 2126
rect 2833 2074 2850 2126
rect 2700 2070 2850 2074
rect 3080 2126 3230 2130
rect 3080 2074 3097 2126
rect 3149 2074 3161 2126
rect 3213 2074 3230 2126
rect 3080 2070 3230 2074
rect 3460 2126 3610 2130
rect 3460 2074 3477 2126
rect 3529 2074 3541 2126
rect 3593 2074 3610 2126
rect 3460 2070 3610 2074
rect 3840 2126 3990 2130
rect 3840 2074 3857 2126
rect 3909 2074 3921 2126
rect 3973 2074 3990 2126
rect 3840 2070 3990 2074
rect 2500 1376 2580 1390
rect 2500 1324 2514 1376
rect 2566 1324 2580 1376
rect 2500 1286 2580 1324
rect 2500 1234 2514 1286
rect 2566 1234 2580 1286
rect 2500 1196 2580 1234
rect 2500 1144 2514 1196
rect 2566 1144 2580 1196
rect 2500 1106 2580 1144
rect 2500 1054 2514 1106
rect 2566 1054 2580 1106
rect 2500 1016 2580 1054
rect 2500 964 2514 1016
rect 2566 964 2580 1016
rect 2500 926 2580 964
rect 2500 874 2514 926
rect 2566 874 2580 926
rect 2500 860 2580 874
rect 2880 1376 2960 1390
rect 2880 1324 2894 1376
rect 2946 1324 2960 1376
rect 2880 1286 2960 1324
rect 2880 1234 2894 1286
rect 2946 1234 2960 1286
rect 2880 1196 2960 1234
rect 2880 1144 2894 1196
rect 2946 1144 2960 1196
rect 2880 1106 2960 1144
rect 2880 1054 2894 1106
rect 2946 1054 2960 1106
rect 2880 1016 2960 1054
rect 2880 964 2894 1016
rect 2946 964 2960 1016
rect 2880 926 2960 964
rect 2880 874 2894 926
rect 2946 874 2960 926
rect 2880 860 2960 874
rect 3260 1376 3340 1390
rect 3260 1324 3274 1376
rect 3326 1324 3340 1376
rect 3260 1286 3340 1324
rect 3260 1234 3274 1286
rect 3326 1234 3340 1286
rect 3260 1196 3340 1234
rect 3260 1144 3274 1196
rect 3326 1144 3340 1196
rect 3260 1106 3340 1144
rect 3260 1054 3274 1106
rect 3326 1054 3340 1106
rect 3260 1016 3340 1054
rect 3260 964 3274 1016
rect 3326 964 3340 1016
rect 3260 926 3340 964
rect 3260 874 3274 926
rect 3326 874 3340 926
rect 3260 860 3340 874
rect 3640 1376 3720 1390
rect 3640 1324 3654 1376
rect 3706 1324 3720 1376
rect 3640 1286 3720 1324
rect 3640 1234 3654 1286
rect 3706 1234 3720 1286
rect 3640 1196 3720 1234
rect 3640 1144 3654 1196
rect 3706 1144 3720 1196
rect 3640 1106 3720 1144
rect 3640 1054 3654 1106
rect 3706 1054 3720 1106
rect 3640 1016 3720 1054
rect 3640 964 3654 1016
rect 3706 964 3720 1016
rect 3640 926 3720 964
rect 3640 874 3654 926
rect 3706 874 3720 926
rect 3640 860 3720 874
rect 4020 1376 4100 1390
rect 4020 1324 4034 1376
rect 4086 1324 4100 1376
rect 4020 1286 4100 1324
rect 4020 1234 4034 1286
rect 4086 1234 4100 1286
rect 4020 1196 4100 1234
rect 4020 1144 4034 1196
rect 4086 1144 4100 1196
rect 4020 1106 4100 1144
rect 4020 1054 4034 1106
rect 4086 1054 4100 1106
rect 4020 1016 4100 1054
rect 4020 964 4034 1016
rect 4086 964 4100 1016
rect 4020 926 4100 964
rect 4020 874 4034 926
rect 4086 874 4100 926
rect 4020 860 4100 874
rect 4130 70 4190 2190
rect 4220 2136 4390 2150
rect 4220 2084 4234 2136
rect 4286 2084 4324 2136
rect 4376 2130 4390 2136
rect 4510 2130 4570 4250
rect 4780 3526 4860 3540
rect 4780 3474 4794 3526
rect 4846 3474 4860 3526
rect 4780 3436 4860 3474
rect 4780 3384 4794 3436
rect 4846 3384 4860 3436
rect 4780 3346 4860 3384
rect 4780 3294 4794 3346
rect 4846 3294 4860 3346
rect 4780 3256 4860 3294
rect 4780 3204 4794 3256
rect 4846 3204 4860 3256
rect 4780 3166 4860 3204
rect 4780 3114 4794 3166
rect 4846 3114 4860 3166
rect 4780 3076 4860 3114
rect 4780 3024 4794 3076
rect 4846 3024 4860 3076
rect 4780 3010 4860 3024
rect 5160 3526 5240 3540
rect 5160 3474 5174 3526
rect 5226 3474 5240 3526
rect 5160 3436 5240 3474
rect 5160 3384 5174 3436
rect 5226 3384 5240 3436
rect 5160 3346 5240 3384
rect 5160 3294 5174 3346
rect 5226 3294 5240 3346
rect 5160 3256 5240 3294
rect 5160 3204 5174 3256
rect 5226 3204 5240 3256
rect 5160 3166 5240 3204
rect 5160 3114 5174 3166
rect 5226 3114 5240 3166
rect 5160 3076 5240 3114
rect 5160 3024 5174 3076
rect 5226 3024 5240 3076
rect 5160 3010 5240 3024
rect 5540 3526 5620 3540
rect 5540 3474 5554 3526
rect 5606 3474 5620 3526
rect 5540 3436 5620 3474
rect 5540 3384 5554 3436
rect 5606 3384 5620 3436
rect 5540 3346 5620 3384
rect 5540 3294 5554 3346
rect 5606 3294 5620 3346
rect 5540 3256 5620 3294
rect 5540 3204 5554 3256
rect 5606 3204 5620 3256
rect 5540 3166 5620 3204
rect 5540 3114 5554 3166
rect 5606 3114 5620 3166
rect 5540 3076 5620 3114
rect 5540 3024 5554 3076
rect 5606 3024 5620 3076
rect 5540 3010 5620 3024
rect 5920 3526 6000 3540
rect 5920 3474 5934 3526
rect 5986 3474 6000 3526
rect 5920 3436 6000 3474
rect 5920 3384 5934 3436
rect 5986 3384 6000 3436
rect 5920 3346 6000 3384
rect 5920 3294 5934 3346
rect 5986 3294 6000 3346
rect 5920 3256 6000 3294
rect 5920 3204 5934 3256
rect 5986 3204 6000 3256
rect 5920 3166 6000 3204
rect 5920 3114 5934 3166
rect 5986 3114 6000 3166
rect 5920 3076 6000 3114
rect 5920 3024 5934 3076
rect 5986 3024 6000 3076
rect 5920 3010 6000 3024
rect 6300 3526 6380 3540
rect 6300 3474 6314 3526
rect 6366 3474 6380 3526
rect 6300 3436 6380 3474
rect 6300 3384 6314 3436
rect 6366 3384 6380 3436
rect 6300 3346 6380 3384
rect 6300 3294 6314 3346
rect 6366 3294 6380 3346
rect 6300 3256 6380 3294
rect 6300 3204 6314 3256
rect 6366 3204 6380 3256
rect 6300 3166 6380 3204
rect 6300 3114 6314 3166
rect 6366 3114 6380 3166
rect 6300 3076 6380 3114
rect 6300 3024 6314 3076
rect 6366 3024 6380 3076
rect 6300 3010 6380 3024
rect 6680 3526 6760 3540
rect 6680 3474 6694 3526
rect 6746 3474 6760 3526
rect 6680 3436 6760 3474
rect 6680 3384 6694 3436
rect 6746 3384 6760 3436
rect 6680 3346 6760 3384
rect 6680 3294 6694 3346
rect 6746 3294 6760 3346
rect 6680 3256 6760 3294
rect 6680 3204 6694 3256
rect 6746 3204 6760 3256
rect 6680 3166 6760 3204
rect 6680 3114 6694 3166
rect 6746 3114 6760 3166
rect 6680 3076 6760 3114
rect 6680 3024 6694 3076
rect 6746 3024 6760 3076
rect 6680 3010 6760 3024
rect 7060 3526 7140 3540
rect 7060 3474 7074 3526
rect 7126 3474 7140 3526
rect 7060 3436 7140 3474
rect 7060 3384 7074 3436
rect 7126 3384 7140 3436
rect 7060 3346 7140 3384
rect 7060 3294 7074 3346
rect 7126 3294 7140 3346
rect 7060 3256 7140 3294
rect 7060 3204 7074 3256
rect 7126 3204 7140 3256
rect 7060 3166 7140 3204
rect 7060 3114 7074 3166
rect 7126 3114 7140 3166
rect 7060 3076 7140 3114
rect 7060 3024 7074 3076
rect 7126 3024 7140 3076
rect 7060 3010 7140 3024
rect 7440 3526 7520 3540
rect 7440 3474 7454 3526
rect 7506 3474 7520 3526
rect 7440 3436 7520 3474
rect 7440 3384 7454 3436
rect 7506 3384 7520 3436
rect 7440 3346 7520 3384
rect 7440 3294 7454 3346
rect 7506 3294 7520 3346
rect 7440 3256 7520 3294
rect 7440 3204 7454 3256
rect 7506 3204 7520 3256
rect 7440 3166 7520 3204
rect 7440 3114 7454 3166
rect 7506 3114 7520 3166
rect 7440 3076 7520 3114
rect 7440 3024 7454 3076
rect 7506 3024 7520 3076
rect 7440 3010 7520 3024
rect 7820 3526 7900 3540
rect 7820 3474 7834 3526
rect 7886 3474 7900 3526
rect 7820 3436 7900 3474
rect 7820 3384 7834 3436
rect 7886 3384 7900 3436
rect 7820 3346 7900 3384
rect 7820 3294 7834 3346
rect 7886 3294 7900 3346
rect 7820 3256 7900 3294
rect 7820 3204 7834 3256
rect 7886 3204 7900 3256
rect 7820 3166 7900 3204
rect 7820 3114 7834 3166
rect 7886 3114 7900 3166
rect 7820 3076 7900 3114
rect 7820 3024 7834 3076
rect 7886 3024 7900 3076
rect 7820 3010 7900 3024
rect 8200 3526 8280 3540
rect 8200 3474 8214 3526
rect 8266 3474 8280 3526
rect 8200 3436 8280 3474
rect 8200 3384 8214 3436
rect 8266 3384 8280 3436
rect 8200 3346 8280 3384
rect 8200 3294 8214 3346
rect 8266 3294 8280 3346
rect 8200 3256 8280 3294
rect 8200 3204 8214 3256
rect 8266 3204 8280 3256
rect 8200 3166 8280 3204
rect 8200 3114 8214 3166
rect 8266 3114 8280 3166
rect 8200 3076 8280 3114
rect 8200 3024 8214 3076
rect 8266 3024 8280 3076
rect 8200 3010 8280 3024
rect 8600 2250 8660 4250
rect 4600 2246 4750 2250
rect 4600 2194 4617 2246
rect 4669 2194 4681 2246
rect 4733 2194 4750 2246
rect 4600 2190 4750 2194
rect 4980 2246 5130 2250
rect 4980 2194 4997 2246
rect 5049 2194 5061 2246
rect 5113 2194 5130 2246
rect 4980 2190 5130 2194
rect 5360 2246 5510 2250
rect 5360 2194 5377 2246
rect 5429 2194 5441 2246
rect 5493 2194 5510 2246
rect 5360 2190 5510 2194
rect 5740 2246 5890 2250
rect 5740 2194 5757 2246
rect 5809 2194 5821 2246
rect 5873 2194 5890 2246
rect 5740 2190 5890 2194
rect 6120 2246 6270 2250
rect 6120 2194 6137 2246
rect 6189 2194 6201 2246
rect 6253 2194 6270 2246
rect 6120 2190 6270 2194
rect 6500 2246 6650 2250
rect 6500 2194 6517 2246
rect 6569 2194 6581 2246
rect 6633 2194 6650 2246
rect 6500 2190 6650 2194
rect 6880 2246 7030 2250
rect 6880 2194 6897 2246
rect 6949 2194 6961 2246
rect 7013 2194 7030 2246
rect 6880 2190 7030 2194
rect 7260 2246 7410 2250
rect 7260 2194 7277 2246
rect 7329 2194 7341 2246
rect 7393 2194 7410 2246
rect 7260 2190 7410 2194
rect 7640 2246 7790 2250
rect 7640 2194 7657 2246
rect 7709 2194 7721 2246
rect 7773 2194 7790 2246
rect 7640 2190 7790 2194
rect 8020 2246 8170 2250
rect 8020 2194 8037 2246
rect 8089 2194 8101 2246
rect 8153 2194 8170 2246
rect 8020 2190 8170 2194
rect 4376 2084 4480 2130
rect 4220 2070 4480 2084
rect 4510 2126 4750 2130
rect 4510 2074 4617 2126
rect 4669 2074 4681 2126
rect 4733 2074 4750 2126
rect 4510 2070 4750 2074
rect 4980 2126 5130 2130
rect 4980 2074 4997 2126
rect 5049 2074 5061 2126
rect 5113 2074 5130 2126
rect 4980 2070 5130 2074
rect 5360 2126 5510 2130
rect 5360 2074 5377 2126
rect 5429 2074 5441 2126
rect 5493 2074 5510 2126
rect 5360 2070 5510 2074
rect 5740 2126 5890 2130
rect 5740 2074 5757 2126
rect 5809 2074 5821 2126
rect 5873 2074 5890 2126
rect 5740 2070 5890 2074
rect 6120 2126 6270 2130
rect 6120 2074 6137 2126
rect 6189 2074 6201 2126
rect 6253 2074 6270 2126
rect 6120 2070 6270 2074
rect 6500 2126 6650 2130
rect 6500 2074 6517 2126
rect 6569 2074 6581 2126
rect 6633 2074 6650 2126
rect 6500 2070 6650 2074
rect 6880 2126 7030 2130
rect 6880 2074 6897 2126
rect 6949 2074 6961 2126
rect 7013 2074 7030 2126
rect 6880 2070 7030 2074
rect 7260 2126 7410 2130
rect 7260 2074 7277 2126
rect 7329 2074 7341 2126
rect 7393 2074 7410 2126
rect 7260 2070 7410 2074
rect 7640 2126 7790 2130
rect 7640 2074 7657 2126
rect 7709 2074 7721 2126
rect 7773 2074 7790 2126
rect 7640 2070 7790 2074
rect 8020 2126 8170 2130
rect 8020 2074 8037 2126
rect 8089 2074 8101 2126
rect 8153 2074 8170 2126
rect 8020 2070 8170 2074
rect 8370 2070 8660 2250
rect -150 2 300 70
rect 420 66 570 70
rect 420 14 437 66
rect 489 14 501 66
rect 553 14 570 66
rect 420 10 570 14
rect 800 66 950 70
rect 800 14 817 66
rect 869 14 881 66
rect 933 14 950 66
rect 800 10 950 14
rect 1180 66 1330 70
rect 1180 14 1197 66
rect 1249 14 1261 66
rect 1313 14 1330 66
rect 1180 10 1330 14
rect 1560 66 1710 70
rect 1560 14 1577 66
rect 1629 14 1641 66
rect 1693 14 1710 66
rect 1560 10 1710 14
rect 1940 66 2090 70
rect 1940 14 1957 66
rect 2009 14 2021 66
rect 2073 14 2090 66
rect 1940 10 2090 14
rect 2230 66 2470 70
rect 2230 14 2337 66
rect 2389 14 2401 66
rect 2453 14 2470 66
rect 2230 10 2470 14
rect 2700 66 2850 70
rect 2700 14 2717 66
rect 2769 14 2781 66
rect 2833 14 2850 66
rect 2700 10 2850 14
rect 3080 66 3230 70
rect 3080 14 3097 66
rect 3149 14 3161 66
rect 3213 14 3230 66
rect 3080 10 3230 14
rect 3460 66 3610 70
rect 3460 14 3477 66
rect 3529 14 3541 66
rect 3593 14 3610 66
rect 3460 10 3610 14
rect 3840 66 3990 70
rect 3840 14 3857 66
rect 3909 14 3921 66
rect 3973 14 3990 66
rect 3840 10 3990 14
rect 4050 27 4370 70
rect -150 -32 -92 2
rect -58 -32 300 2
rect -150 -110 300 -32
rect 4050 -7 4093 27
rect 4127 10 4370 27
rect 4127 -7 4190 10
rect 4050 -50 4190 -7
rect 4420 -50 4480 2070
rect 4780 1376 4860 1390
rect 4780 1324 4794 1376
rect 4846 1324 4860 1376
rect 4780 1286 4860 1324
rect 4780 1234 4794 1286
rect 4846 1234 4860 1286
rect 4780 1196 4860 1234
rect 4780 1144 4794 1196
rect 4846 1144 4860 1196
rect 4780 1106 4860 1144
rect 4780 1054 4794 1106
rect 4846 1054 4860 1106
rect 4780 1016 4860 1054
rect 4780 964 4794 1016
rect 4846 964 4860 1016
rect 4780 926 4860 964
rect 4780 874 4794 926
rect 4846 874 4860 926
rect 4780 860 4860 874
rect 5160 1376 5240 1390
rect 5160 1324 5174 1376
rect 5226 1324 5240 1376
rect 5160 1286 5240 1324
rect 5160 1234 5174 1286
rect 5226 1234 5240 1286
rect 5160 1196 5240 1234
rect 5160 1144 5174 1196
rect 5226 1144 5240 1196
rect 5160 1106 5240 1144
rect 5160 1054 5174 1106
rect 5226 1054 5240 1106
rect 5160 1016 5240 1054
rect 5160 964 5174 1016
rect 5226 964 5240 1016
rect 5160 926 5240 964
rect 5160 874 5174 926
rect 5226 874 5240 926
rect 5160 860 5240 874
rect 5540 1376 5620 1390
rect 5540 1324 5554 1376
rect 5606 1324 5620 1376
rect 5540 1286 5620 1324
rect 5540 1234 5554 1286
rect 5606 1234 5620 1286
rect 5540 1196 5620 1234
rect 5540 1144 5554 1196
rect 5606 1144 5620 1196
rect 5540 1106 5620 1144
rect 5540 1054 5554 1106
rect 5606 1054 5620 1106
rect 5540 1016 5620 1054
rect 5540 964 5554 1016
rect 5606 964 5620 1016
rect 5540 926 5620 964
rect 5540 874 5554 926
rect 5606 874 5620 926
rect 5540 860 5620 874
rect 5920 1376 6000 1390
rect 5920 1324 5934 1376
rect 5986 1324 6000 1376
rect 5920 1286 6000 1324
rect 5920 1234 5934 1286
rect 5986 1234 6000 1286
rect 5920 1196 6000 1234
rect 5920 1144 5934 1196
rect 5986 1144 6000 1196
rect 5920 1106 6000 1144
rect 5920 1054 5934 1106
rect 5986 1054 6000 1106
rect 5920 1016 6000 1054
rect 5920 964 5934 1016
rect 5986 964 6000 1016
rect 5920 926 6000 964
rect 5920 874 5934 926
rect 5986 874 6000 926
rect 5920 860 6000 874
rect 6300 1376 6380 1390
rect 6300 1324 6314 1376
rect 6366 1324 6380 1376
rect 6300 1286 6380 1324
rect 6300 1234 6314 1286
rect 6366 1234 6380 1286
rect 6300 1196 6380 1234
rect 6300 1144 6314 1196
rect 6366 1144 6380 1196
rect 6300 1106 6380 1144
rect 6300 1054 6314 1106
rect 6366 1054 6380 1106
rect 6300 1016 6380 1054
rect 6300 964 6314 1016
rect 6366 964 6380 1016
rect 6300 926 6380 964
rect 6300 874 6314 926
rect 6366 874 6380 926
rect 6300 860 6380 874
rect 6680 1376 6760 1390
rect 6680 1324 6694 1376
rect 6746 1324 6760 1376
rect 6680 1286 6760 1324
rect 6680 1234 6694 1286
rect 6746 1234 6760 1286
rect 6680 1196 6760 1234
rect 6680 1144 6694 1196
rect 6746 1144 6760 1196
rect 6680 1106 6760 1144
rect 6680 1054 6694 1106
rect 6746 1054 6760 1106
rect 6680 1016 6760 1054
rect 6680 964 6694 1016
rect 6746 964 6760 1016
rect 6680 926 6760 964
rect 6680 874 6694 926
rect 6746 874 6760 926
rect 6680 860 6760 874
rect 7060 1376 7140 1390
rect 7060 1324 7074 1376
rect 7126 1324 7140 1376
rect 7060 1286 7140 1324
rect 7060 1234 7074 1286
rect 7126 1234 7140 1286
rect 7060 1196 7140 1234
rect 7060 1144 7074 1196
rect 7126 1144 7140 1196
rect 7060 1106 7140 1144
rect 7060 1054 7074 1106
rect 7126 1054 7140 1106
rect 7060 1016 7140 1054
rect 7060 964 7074 1016
rect 7126 964 7140 1016
rect 7060 926 7140 964
rect 7060 874 7074 926
rect 7126 874 7140 926
rect 7060 860 7140 874
rect 7440 1376 7520 1390
rect 7440 1324 7454 1376
rect 7506 1324 7520 1376
rect 7440 1286 7520 1324
rect 7440 1234 7454 1286
rect 7506 1234 7520 1286
rect 7440 1196 7520 1234
rect 7440 1144 7454 1196
rect 7506 1144 7520 1196
rect 7440 1106 7520 1144
rect 7440 1054 7454 1106
rect 7506 1054 7520 1106
rect 7440 1016 7520 1054
rect 7440 964 7454 1016
rect 7506 964 7520 1016
rect 7440 926 7520 964
rect 7440 874 7454 926
rect 7506 874 7520 926
rect 7440 860 7520 874
rect 7820 1376 7900 1390
rect 7820 1324 7834 1376
rect 7886 1324 7900 1376
rect 7820 1286 7900 1324
rect 7820 1234 7834 1286
rect 7886 1234 7900 1286
rect 7820 1196 7900 1234
rect 7820 1144 7834 1196
rect 7886 1144 7900 1196
rect 7820 1106 7900 1144
rect 7820 1054 7834 1106
rect 7886 1054 7900 1106
rect 7820 1016 7900 1054
rect 7820 964 7834 1016
rect 7886 964 7900 1016
rect 7820 926 7900 964
rect 7820 874 7834 926
rect 7886 874 7900 926
rect 7820 860 7900 874
rect 8200 1376 8280 1390
rect 8200 1324 8214 1376
rect 8266 1324 8280 1376
rect 8200 1286 8280 1324
rect 8200 1234 8214 1286
rect 8266 1234 8280 1286
rect 8200 1196 8280 1234
rect 8200 1144 8214 1196
rect 8266 1144 8280 1196
rect 8200 1106 8280 1144
rect 8200 1054 8214 1106
rect 8266 1054 8280 1106
rect 8200 1016 8280 1054
rect 8200 964 8214 1016
rect 8266 964 8280 1016
rect 8200 926 8280 964
rect 8200 874 8214 926
rect 8266 874 8280 926
rect 8200 860 8280 874
rect 8600 70 8660 2070
rect 8830 4306 8910 5020
rect 8830 4254 8844 4306
rect 8896 4254 8910 4306
rect 8830 4226 8910 4254
rect 8830 4174 8844 4226
rect 8896 4174 8910 4226
rect 8830 2126 8910 4174
rect 8830 2074 8844 2126
rect 8896 2074 8910 2126
rect 8830 2046 8910 2074
rect 8830 1994 8844 2046
rect 8896 1994 8910 2046
rect 8830 1990 8910 1994
rect 4600 66 4750 70
rect 4600 14 4617 66
rect 4669 14 4681 66
rect 4733 14 4750 66
rect 4600 10 4750 14
rect 4980 66 5130 70
rect 4980 14 4997 66
rect 5049 14 5061 66
rect 5113 14 5130 66
rect 4980 10 5130 14
rect 5360 66 5510 70
rect 5360 14 5377 66
rect 5429 14 5441 66
rect 5493 14 5510 66
rect 5360 10 5510 14
rect 5740 66 5890 70
rect 5740 14 5757 66
rect 5809 14 5821 66
rect 5873 14 5890 66
rect 5740 10 5890 14
rect 6120 66 6270 70
rect 6120 14 6137 66
rect 6189 14 6201 66
rect 6253 14 6270 66
rect 6120 10 6270 14
rect 6500 66 6650 70
rect 6500 14 6517 66
rect 6569 14 6581 66
rect 6633 14 6650 66
rect 6500 10 6650 14
rect 6880 66 7030 70
rect 6880 14 6897 66
rect 6949 14 6961 66
rect 7013 14 7030 66
rect 6880 10 7030 14
rect 7260 66 7410 70
rect 7260 14 7277 66
rect 7329 14 7341 66
rect 7393 14 7410 66
rect 7260 10 7410 14
rect 7640 66 7790 70
rect 7640 14 7657 66
rect 7709 14 7721 66
rect 7773 14 7790 66
rect 7640 10 7790 14
rect 8020 66 8170 70
rect 8020 14 8037 66
rect 8089 14 8101 66
rect 8153 14 8170 66
rect 8020 10 8170 14
rect 420 -54 570 -50
rect 420 -106 437 -54
rect 489 -106 501 -54
rect 553 -106 570 -54
rect 420 -110 570 -106
rect 800 -54 950 -50
rect 800 -106 817 -54
rect 869 -106 881 -54
rect 933 -106 950 -54
rect 800 -110 950 -106
rect 1180 -54 1330 -50
rect 1180 -106 1197 -54
rect 1249 -106 1261 -54
rect 1313 -106 1330 -54
rect 1180 -110 1330 -106
rect 1560 -54 1710 -50
rect 1560 -106 1577 -54
rect 1629 -106 1641 -54
rect 1693 -106 1710 -54
rect 1560 -110 1710 -106
rect 1940 -54 2090 -50
rect 1940 -106 1957 -54
rect 2009 -106 2021 -54
rect 2073 -106 2090 -54
rect 1940 -110 2090 -106
rect 2320 -54 2470 -50
rect 2320 -106 2337 -54
rect 2389 -106 2401 -54
rect 2453 -106 2470 -54
rect 2320 -110 2470 -106
rect 2700 -54 2850 -50
rect 2700 -106 2717 -54
rect 2769 -106 2781 -54
rect 2833 -106 2850 -54
rect 2700 -110 2850 -106
rect 3080 -54 3230 -50
rect 3080 -106 3097 -54
rect 3149 -106 3161 -54
rect 3213 -106 3230 -54
rect 3080 -110 3230 -106
rect 3460 -54 3610 -50
rect 3460 -106 3477 -54
rect 3529 -106 3541 -54
rect 3593 -106 3610 -54
rect 3460 -110 3610 -106
rect 3840 -54 3990 -50
rect 3840 -106 3857 -54
rect 3909 -106 3921 -54
rect 3973 -106 3990 -54
rect 3840 -110 3990 -106
rect 4220 -110 4480 -50
rect 4600 -54 4750 -50
rect 4600 -106 4617 -54
rect 4669 -106 4681 -54
rect 4733 -106 4750 -54
rect 4600 -110 4750 -106
rect 4980 -54 5130 -50
rect 4980 -106 4997 -54
rect 5049 -106 5061 -54
rect 5113 -106 5130 -54
rect 4980 -110 5130 -106
rect 5360 -54 5510 -50
rect 5360 -106 5377 -54
rect 5429 -106 5441 -54
rect 5493 -106 5510 -54
rect 5360 -110 5510 -106
rect 5740 -54 5890 -50
rect 5740 -106 5757 -54
rect 5809 -106 5821 -54
rect 5873 -106 5890 -54
rect 5740 -110 5890 -106
rect 6120 -54 6270 -50
rect 6120 -106 6137 -54
rect 6189 -106 6201 -54
rect 6253 -106 6270 -54
rect 6120 -110 6270 -106
rect 6500 -54 6650 -50
rect 6500 -106 6517 -54
rect 6569 -106 6581 -54
rect 6633 -106 6650 -54
rect 6500 -110 6650 -106
rect 6880 -54 7030 -50
rect 6880 -106 6897 -54
rect 6949 -106 6961 -54
rect 7013 -106 7030 -54
rect 6880 -110 7030 -106
rect 7260 -54 7410 -50
rect 7260 -106 7277 -54
rect 7329 -106 7341 -54
rect 7393 -106 7410 -54
rect 7260 -110 7410 -106
rect 7640 -54 7790 -50
rect 7640 -106 7657 -54
rect 7709 -106 7721 -54
rect 7773 -106 7790 -54
rect 7640 -110 7790 -106
rect 8020 -54 8170 -50
rect 8020 -106 8037 -54
rect 8089 -106 8101 -54
rect 8153 -106 8170 -54
rect 8020 -110 8170 -106
rect 8370 -110 8660 70
rect -250 -2034 -170 -2030
rect -250 -2086 -236 -2034
rect -184 -2086 -170 -2034
rect -250 -2114 -170 -2086
rect 240 -2110 300 -110
rect 600 -864 680 -850
rect 600 -916 614 -864
rect 666 -916 680 -864
rect 600 -954 680 -916
rect 600 -1006 614 -954
rect 666 -1006 680 -954
rect 600 -1044 680 -1006
rect 600 -1096 614 -1044
rect 666 -1096 680 -1044
rect 600 -1134 680 -1096
rect 600 -1186 614 -1134
rect 666 -1186 680 -1134
rect 600 -1224 680 -1186
rect 600 -1276 614 -1224
rect 666 -1276 680 -1224
rect 600 -1314 680 -1276
rect 600 -1366 614 -1314
rect 666 -1366 680 -1314
rect 600 -1380 680 -1366
rect 980 -864 1060 -850
rect 980 -916 994 -864
rect 1046 -916 1060 -864
rect 980 -954 1060 -916
rect 980 -1006 994 -954
rect 1046 -1006 1060 -954
rect 980 -1044 1060 -1006
rect 980 -1096 994 -1044
rect 1046 -1096 1060 -1044
rect 980 -1134 1060 -1096
rect 980 -1186 994 -1134
rect 1046 -1186 1060 -1134
rect 980 -1224 1060 -1186
rect 980 -1276 994 -1224
rect 1046 -1276 1060 -1224
rect 980 -1314 1060 -1276
rect 980 -1366 994 -1314
rect 1046 -1366 1060 -1314
rect 980 -1380 1060 -1366
rect 1360 -864 1440 -850
rect 1360 -916 1374 -864
rect 1426 -916 1440 -864
rect 1360 -954 1440 -916
rect 1360 -1006 1374 -954
rect 1426 -1006 1440 -954
rect 1360 -1044 1440 -1006
rect 1360 -1096 1374 -1044
rect 1426 -1096 1440 -1044
rect 1360 -1134 1440 -1096
rect 1360 -1186 1374 -1134
rect 1426 -1186 1440 -1134
rect 1360 -1224 1440 -1186
rect 1360 -1276 1374 -1224
rect 1426 -1276 1440 -1224
rect 1360 -1314 1440 -1276
rect 1360 -1366 1374 -1314
rect 1426 -1366 1440 -1314
rect 1360 -1380 1440 -1366
rect 1740 -864 1820 -850
rect 1740 -916 1754 -864
rect 1806 -916 1820 -864
rect 1740 -954 1820 -916
rect 1740 -1006 1754 -954
rect 1806 -1006 1820 -954
rect 1740 -1044 1820 -1006
rect 1740 -1096 1754 -1044
rect 1806 -1096 1820 -1044
rect 1740 -1134 1820 -1096
rect 1740 -1186 1754 -1134
rect 1806 -1186 1820 -1134
rect 1740 -1224 1820 -1186
rect 1740 -1276 1754 -1224
rect 1806 -1276 1820 -1224
rect 1740 -1314 1820 -1276
rect 1740 -1366 1754 -1314
rect 1806 -1366 1820 -1314
rect 1740 -1380 1820 -1366
rect 2120 -864 2200 -850
rect 2120 -916 2134 -864
rect 2186 -916 2200 -864
rect 2120 -954 2200 -916
rect 2120 -1006 2134 -954
rect 2186 -1006 2200 -954
rect 2120 -1044 2200 -1006
rect 2120 -1096 2134 -1044
rect 2186 -1096 2200 -1044
rect 2120 -1134 2200 -1096
rect 2120 -1186 2134 -1134
rect 2186 -1186 2200 -1134
rect 2120 -1224 2200 -1186
rect 2120 -1276 2134 -1224
rect 2186 -1276 2200 -1224
rect 2120 -1314 2200 -1276
rect 2120 -1366 2134 -1314
rect 2186 -1366 2200 -1314
rect 2120 -1380 2200 -1366
rect 2500 -864 2580 -850
rect 2500 -916 2514 -864
rect 2566 -916 2580 -864
rect 2500 -954 2580 -916
rect 2500 -1006 2514 -954
rect 2566 -1006 2580 -954
rect 2500 -1044 2580 -1006
rect 2500 -1096 2514 -1044
rect 2566 -1096 2580 -1044
rect 2500 -1134 2580 -1096
rect 2500 -1186 2514 -1134
rect 2566 -1186 2580 -1134
rect 2500 -1224 2580 -1186
rect 2500 -1276 2514 -1224
rect 2566 -1276 2580 -1224
rect 2500 -1314 2580 -1276
rect 2500 -1366 2514 -1314
rect 2566 -1366 2580 -1314
rect 2500 -1380 2580 -1366
rect 2880 -864 2960 -850
rect 2880 -916 2894 -864
rect 2946 -916 2960 -864
rect 2880 -954 2960 -916
rect 2880 -1006 2894 -954
rect 2946 -1006 2960 -954
rect 2880 -1044 2960 -1006
rect 2880 -1096 2894 -1044
rect 2946 -1096 2960 -1044
rect 2880 -1134 2960 -1096
rect 2880 -1186 2894 -1134
rect 2946 -1186 2960 -1134
rect 2880 -1224 2960 -1186
rect 2880 -1276 2894 -1224
rect 2946 -1276 2960 -1224
rect 2880 -1314 2960 -1276
rect 2880 -1366 2894 -1314
rect 2946 -1366 2960 -1314
rect 2880 -1380 2960 -1366
rect 3260 -864 3340 -850
rect 3260 -916 3274 -864
rect 3326 -916 3340 -864
rect 3260 -954 3340 -916
rect 3260 -1006 3274 -954
rect 3326 -1006 3340 -954
rect 3260 -1044 3340 -1006
rect 3260 -1096 3274 -1044
rect 3326 -1096 3340 -1044
rect 3260 -1134 3340 -1096
rect 3260 -1186 3274 -1134
rect 3326 -1186 3340 -1134
rect 3260 -1224 3340 -1186
rect 3260 -1276 3274 -1224
rect 3326 -1276 3340 -1224
rect 3260 -1314 3340 -1276
rect 3260 -1366 3274 -1314
rect 3326 -1366 3340 -1314
rect 3260 -1380 3340 -1366
rect 3640 -864 3720 -850
rect 3640 -916 3654 -864
rect 3706 -916 3720 -864
rect 3640 -954 3720 -916
rect 3640 -1006 3654 -954
rect 3706 -1006 3720 -954
rect 3640 -1044 3720 -1006
rect 3640 -1096 3654 -1044
rect 3706 -1096 3720 -1044
rect 3640 -1134 3720 -1096
rect 3640 -1186 3654 -1134
rect 3706 -1186 3720 -1134
rect 3640 -1224 3720 -1186
rect 3640 -1276 3654 -1224
rect 3706 -1276 3720 -1224
rect 3640 -1314 3720 -1276
rect 3640 -1366 3654 -1314
rect 3706 -1366 3720 -1314
rect 3640 -1380 3720 -1366
rect 4020 -864 4100 -850
rect 4020 -916 4034 -864
rect 4086 -916 4100 -864
rect 4020 -954 4100 -916
rect 4020 -1006 4034 -954
rect 4086 -1006 4100 -954
rect 4020 -1044 4100 -1006
rect 4020 -1096 4034 -1044
rect 4086 -1096 4100 -1044
rect 4020 -1134 4100 -1096
rect 4020 -1186 4034 -1134
rect 4086 -1186 4100 -1134
rect 4020 -1224 4100 -1186
rect 4020 -1276 4034 -1224
rect 4086 -1276 4100 -1224
rect 4020 -1314 4100 -1276
rect 4020 -1366 4034 -1314
rect 4086 -1366 4100 -1314
rect 4020 -1380 4100 -1366
rect 4420 -1820 4480 -110
rect 4780 -864 4860 -850
rect 4780 -916 4794 -864
rect 4846 -916 4860 -864
rect 4780 -954 4860 -916
rect 4780 -1006 4794 -954
rect 4846 -1006 4860 -954
rect 4780 -1044 4860 -1006
rect 4780 -1096 4794 -1044
rect 4846 -1096 4860 -1044
rect 4780 -1134 4860 -1096
rect 4780 -1186 4794 -1134
rect 4846 -1186 4860 -1134
rect 4780 -1224 4860 -1186
rect 4780 -1276 4794 -1224
rect 4846 -1276 4860 -1224
rect 4780 -1314 4860 -1276
rect 4780 -1366 4794 -1314
rect 4846 -1366 4860 -1314
rect 4780 -1380 4860 -1366
rect 5160 -864 5240 -850
rect 5160 -916 5174 -864
rect 5226 -916 5240 -864
rect 5160 -954 5240 -916
rect 5160 -1006 5174 -954
rect 5226 -1006 5240 -954
rect 5160 -1044 5240 -1006
rect 5160 -1096 5174 -1044
rect 5226 -1096 5240 -1044
rect 5160 -1134 5240 -1096
rect 5160 -1186 5174 -1134
rect 5226 -1186 5240 -1134
rect 5160 -1224 5240 -1186
rect 5160 -1276 5174 -1224
rect 5226 -1276 5240 -1224
rect 5160 -1314 5240 -1276
rect 5160 -1366 5174 -1314
rect 5226 -1366 5240 -1314
rect 5160 -1380 5240 -1366
rect 5540 -864 5620 -850
rect 5540 -916 5554 -864
rect 5606 -916 5620 -864
rect 5540 -954 5620 -916
rect 5540 -1006 5554 -954
rect 5606 -1006 5620 -954
rect 5540 -1044 5620 -1006
rect 5540 -1096 5554 -1044
rect 5606 -1096 5620 -1044
rect 5540 -1134 5620 -1096
rect 5540 -1186 5554 -1134
rect 5606 -1186 5620 -1134
rect 5540 -1224 5620 -1186
rect 5540 -1276 5554 -1224
rect 5606 -1276 5620 -1224
rect 5540 -1314 5620 -1276
rect 5540 -1366 5554 -1314
rect 5606 -1366 5620 -1314
rect 5540 -1380 5620 -1366
rect 5920 -864 6000 -850
rect 5920 -916 5934 -864
rect 5986 -916 6000 -864
rect 5920 -954 6000 -916
rect 5920 -1006 5934 -954
rect 5986 -1006 6000 -954
rect 5920 -1044 6000 -1006
rect 5920 -1096 5934 -1044
rect 5986 -1096 6000 -1044
rect 5920 -1134 6000 -1096
rect 5920 -1186 5934 -1134
rect 5986 -1186 6000 -1134
rect 5920 -1224 6000 -1186
rect 5920 -1276 5934 -1224
rect 5986 -1276 6000 -1224
rect 5920 -1314 6000 -1276
rect 5920 -1366 5934 -1314
rect 5986 -1366 6000 -1314
rect 5920 -1380 6000 -1366
rect 6300 -864 6380 -850
rect 6300 -916 6314 -864
rect 6366 -916 6380 -864
rect 6300 -954 6380 -916
rect 6300 -1006 6314 -954
rect 6366 -1006 6380 -954
rect 6300 -1044 6380 -1006
rect 6300 -1096 6314 -1044
rect 6366 -1096 6380 -1044
rect 6300 -1134 6380 -1096
rect 6300 -1186 6314 -1134
rect 6366 -1186 6380 -1134
rect 6300 -1224 6380 -1186
rect 6300 -1276 6314 -1224
rect 6366 -1276 6380 -1224
rect 6300 -1314 6380 -1276
rect 6300 -1366 6314 -1314
rect 6366 -1366 6380 -1314
rect 6300 -1380 6380 -1366
rect 6680 -864 6760 -850
rect 6680 -916 6694 -864
rect 6746 -916 6760 -864
rect 6680 -954 6760 -916
rect 6680 -1006 6694 -954
rect 6746 -1006 6760 -954
rect 6680 -1044 6760 -1006
rect 6680 -1096 6694 -1044
rect 6746 -1096 6760 -1044
rect 6680 -1134 6760 -1096
rect 6680 -1186 6694 -1134
rect 6746 -1186 6760 -1134
rect 6680 -1224 6760 -1186
rect 6680 -1276 6694 -1224
rect 6746 -1276 6760 -1224
rect 6680 -1314 6760 -1276
rect 6680 -1366 6694 -1314
rect 6746 -1366 6760 -1314
rect 6680 -1380 6760 -1366
rect 7060 -864 7140 -850
rect 7060 -916 7074 -864
rect 7126 -916 7140 -864
rect 7060 -954 7140 -916
rect 7060 -1006 7074 -954
rect 7126 -1006 7140 -954
rect 7060 -1044 7140 -1006
rect 7060 -1096 7074 -1044
rect 7126 -1096 7140 -1044
rect 7060 -1134 7140 -1096
rect 7060 -1186 7074 -1134
rect 7126 -1186 7140 -1134
rect 7060 -1224 7140 -1186
rect 7060 -1276 7074 -1224
rect 7126 -1276 7140 -1224
rect 7060 -1314 7140 -1276
rect 7060 -1366 7074 -1314
rect 7126 -1366 7140 -1314
rect 7060 -1380 7140 -1366
rect 7440 -864 7520 -850
rect 7440 -916 7454 -864
rect 7506 -916 7520 -864
rect 7440 -954 7520 -916
rect 7440 -1006 7454 -954
rect 7506 -1006 7520 -954
rect 7440 -1044 7520 -1006
rect 7440 -1096 7454 -1044
rect 7506 -1096 7520 -1044
rect 7440 -1134 7520 -1096
rect 7440 -1186 7454 -1134
rect 7506 -1186 7520 -1134
rect 7440 -1224 7520 -1186
rect 7440 -1276 7454 -1224
rect 7506 -1276 7520 -1224
rect 7440 -1314 7520 -1276
rect 7440 -1366 7454 -1314
rect 7506 -1366 7520 -1314
rect 7440 -1380 7520 -1366
rect 7820 -864 7900 -850
rect 7820 -916 7834 -864
rect 7886 -916 7900 -864
rect 7820 -954 7900 -916
rect 7820 -1006 7834 -954
rect 7886 -1006 7900 -954
rect 7820 -1044 7900 -1006
rect 7820 -1096 7834 -1044
rect 7886 -1096 7900 -1044
rect 7820 -1134 7900 -1096
rect 7820 -1186 7834 -1134
rect 7886 -1186 7900 -1134
rect 7820 -1224 7900 -1186
rect 7820 -1276 7834 -1224
rect 7886 -1276 7900 -1224
rect 7820 -1314 7900 -1276
rect 7820 -1366 7834 -1314
rect 7886 -1366 7900 -1314
rect 7820 -1380 7900 -1366
rect 8200 -864 8280 -850
rect 8200 -916 8214 -864
rect 8266 -916 8280 -864
rect 8200 -954 8280 -916
rect 8200 -1006 8214 -954
rect 8266 -1006 8280 -954
rect 8200 -1044 8280 -1006
rect 8200 -1096 8214 -1044
rect 8266 -1096 8280 -1044
rect 8200 -1134 8280 -1096
rect 8200 -1186 8214 -1134
rect 8266 -1186 8280 -1134
rect 8200 -1224 8280 -1186
rect 8200 -1276 8214 -1224
rect 8266 -1276 8280 -1224
rect 8200 -1314 8280 -1276
rect 8200 -1366 8214 -1314
rect 8266 -1366 8280 -1314
rect 8200 -1380 8280 -1366
rect 8600 -2110 8660 -110
rect -250 -2166 -236 -2114
rect -184 -2166 -170 -2114
rect -250 -4214 -170 -2166
rect 10 -2290 300 -2110
rect 420 -2114 570 -2110
rect 420 -2166 437 -2114
rect 489 -2166 501 -2114
rect 553 -2166 570 -2114
rect 420 -2170 570 -2166
rect 800 -2114 950 -2110
rect 800 -2166 817 -2114
rect 869 -2166 881 -2114
rect 933 -2166 950 -2114
rect 800 -2170 950 -2166
rect 1180 -2114 1330 -2110
rect 1180 -2166 1197 -2114
rect 1249 -2166 1261 -2114
rect 1313 -2166 1330 -2114
rect 1180 -2170 1330 -2166
rect 1560 -2114 1710 -2110
rect 1560 -2166 1577 -2114
rect 1629 -2166 1641 -2114
rect 1693 -2166 1710 -2114
rect 1560 -2170 1710 -2166
rect 1940 -2114 2090 -2110
rect 1940 -2166 1957 -2114
rect 2009 -2166 2021 -2114
rect 2073 -2166 2090 -2114
rect 1940 -2170 2090 -2166
rect 2320 -2114 2470 -2110
rect 2320 -2166 2337 -2114
rect 2389 -2166 2401 -2114
rect 2453 -2166 2470 -2114
rect 2320 -2170 2470 -2166
rect 2700 -2114 2850 -2110
rect 2700 -2166 2717 -2114
rect 2769 -2166 2781 -2114
rect 2833 -2166 2850 -2114
rect 2700 -2170 2850 -2166
rect 3080 -2114 3230 -2110
rect 3080 -2166 3097 -2114
rect 3149 -2166 3161 -2114
rect 3213 -2166 3230 -2114
rect 3080 -2170 3230 -2166
rect 3460 -2114 3610 -2110
rect 3460 -2166 3477 -2114
rect 3529 -2166 3541 -2114
rect 3593 -2166 3610 -2114
rect 3460 -2170 3610 -2166
rect 3840 -2114 4190 -2110
rect 3840 -2166 3857 -2114
rect 3909 -2166 3921 -2114
rect 3973 -2166 4004 -2114
rect 4056 -2166 4190 -2114
rect 3840 -2170 4190 -2166
rect 420 -2234 570 -2230
rect 420 -2286 437 -2234
rect 489 -2286 501 -2234
rect 553 -2286 570 -2234
rect 420 -2290 570 -2286
rect 800 -2234 950 -2230
rect 800 -2286 817 -2234
rect 869 -2286 881 -2234
rect 933 -2286 950 -2234
rect 800 -2290 950 -2286
rect 1180 -2234 1330 -2230
rect 1180 -2286 1197 -2234
rect 1249 -2286 1261 -2234
rect 1313 -2286 1330 -2234
rect 1180 -2290 1330 -2286
rect 1560 -2234 1710 -2230
rect 1560 -2286 1577 -2234
rect 1629 -2286 1641 -2234
rect 1693 -2286 1710 -2234
rect 1560 -2290 1710 -2286
rect 1940 -2234 2090 -2230
rect 1940 -2286 1957 -2234
rect 2009 -2286 2021 -2234
rect 2073 -2286 2090 -2234
rect 1940 -2290 2090 -2286
rect 2320 -2234 2470 -2230
rect 2320 -2286 2337 -2234
rect 2389 -2286 2401 -2234
rect 2453 -2286 2470 -2234
rect 2320 -2290 2470 -2286
rect 2700 -2234 2850 -2230
rect 2700 -2286 2717 -2234
rect 2769 -2286 2781 -2234
rect 2833 -2286 2850 -2234
rect 2700 -2290 2850 -2286
rect 3080 -2234 3230 -2230
rect 3080 -2286 3097 -2234
rect 3149 -2286 3161 -2234
rect 3213 -2286 3230 -2234
rect 3080 -2290 3230 -2286
rect 3460 -2234 3610 -2230
rect 3460 -2286 3477 -2234
rect 3529 -2286 3541 -2234
rect 3593 -2286 3610 -2234
rect 3460 -2290 3610 -2286
rect 3840 -2234 3990 -2230
rect 3840 -2286 3857 -2234
rect 3909 -2286 3921 -2234
rect 3973 -2286 3990 -2234
rect 3840 -2290 3990 -2286
rect -250 -4266 -236 -4214
rect -184 -4266 -170 -4214
rect -250 -4294 -170 -4266
rect 220 -4290 300 -2290
rect 600 -3054 680 -3040
rect 600 -3106 614 -3054
rect 666 -3106 680 -3054
rect 600 -3144 680 -3106
rect 600 -3196 614 -3144
rect 666 -3196 680 -3144
rect 600 -3234 680 -3196
rect 600 -3286 614 -3234
rect 666 -3286 680 -3234
rect 600 -3324 680 -3286
rect 600 -3376 614 -3324
rect 666 -3376 680 -3324
rect 600 -3414 680 -3376
rect 600 -3466 614 -3414
rect 666 -3466 680 -3414
rect 600 -3504 680 -3466
rect 600 -3556 614 -3504
rect 666 -3556 680 -3504
rect 600 -3570 680 -3556
rect 980 -3054 1060 -3040
rect 980 -3106 994 -3054
rect 1046 -3106 1060 -3054
rect 980 -3144 1060 -3106
rect 980 -3196 994 -3144
rect 1046 -3196 1060 -3144
rect 980 -3234 1060 -3196
rect 980 -3286 994 -3234
rect 1046 -3286 1060 -3234
rect 980 -3324 1060 -3286
rect 980 -3376 994 -3324
rect 1046 -3376 1060 -3324
rect 980 -3414 1060 -3376
rect 980 -3466 994 -3414
rect 1046 -3466 1060 -3414
rect 980 -3504 1060 -3466
rect 980 -3556 994 -3504
rect 1046 -3556 1060 -3504
rect 980 -3570 1060 -3556
rect 1360 -3054 1440 -3040
rect 1360 -3106 1374 -3054
rect 1426 -3106 1440 -3054
rect 1360 -3144 1440 -3106
rect 1360 -3196 1374 -3144
rect 1426 -3196 1440 -3144
rect 1360 -3234 1440 -3196
rect 1360 -3286 1374 -3234
rect 1426 -3286 1440 -3234
rect 1360 -3324 1440 -3286
rect 1360 -3376 1374 -3324
rect 1426 -3376 1440 -3324
rect 1360 -3414 1440 -3376
rect 1360 -3466 1374 -3414
rect 1426 -3466 1440 -3414
rect 1360 -3504 1440 -3466
rect 1360 -3556 1374 -3504
rect 1426 -3556 1440 -3504
rect 1360 -3570 1440 -3556
rect 1740 -3054 1820 -3040
rect 1740 -3106 1754 -3054
rect 1806 -3106 1820 -3054
rect 1740 -3144 1820 -3106
rect 1740 -3196 1754 -3144
rect 1806 -3196 1820 -3144
rect 1740 -3234 1820 -3196
rect 1740 -3286 1754 -3234
rect 1806 -3286 1820 -3234
rect 1740 -3324 1820 -3286
rect 1740 -3376 1754 -3324
rect 1806 -3376 1820 -3324
rect 1740 -3414 1820 -3376
rect 1740 -3466 1754 -3414
rect 1806 -3466 1820 -3414
rect 1740 -3504 1820 -3466
rect 1740 -3556 1754 -3504
rect 1806 -3556 1820 -3504
rect 1740 -3570 1820 -3556
rect 2120 -3054 2200 -3040
rect 2120 -3106 2134 -3054
rect 2186 -3106 2200 -3054
rect 2120 -3144 2200 -3106
rect 2120 -3196 2134 -3144
rect 2186 -3196 2200 -3144
rect 2120 -3234 2200 -3196
rect 2120 -3286 2134 -3234
rect 2186 -3286 2200 -3234
rect 2120 -3324 2200 -3286
rect 2120 -3376 2134 -3324
rect 2186 -3376 2200 -3324
rect 2120 -3414 2200 -3376
rect 2120 -3466 2134 -3414
rect 2186 -3466 2200 -3414
rect 2120 -3504 2200 -3466
rect 2120 -3556 2134 -3504
rect 2186 -3556 2200 -3504
rect 2120 -3570 2200 -3556
rect 2500 -3054 2580 -3040
rect 2500 -3106 2514 -3054
rect 2566 -3106 2580 -3054
rect 2500 -3144 2580 -3106
rect 2500 -3196 2514 -3144
rect 2566 -3196 2580 -3144
rect 2500 -3234 2580 -3196
rect 2500 -3286 2514 -3234
rect 2566 -3286 2580 -3234
rect 2500 -3324 2580 -3286
rect 2500 -3376 2514 -3324
rect 2566 -3376 2580 -3324
rect 2500 -3414 2580 -3376
rect 2500 -3466 2514 -3414
rect 2566 -3466 2580 -3414
rect 2500 -3504 2580 -3466
rect 2500 -3556 2514 -3504
rect 2566 -3556 2580 -3504
rect 2500 -3570 2580 -3556
rect 2880 -3054 2960 -3040
rect 2880 -3106 2894 -3054
rect 2946 -3106 2960 -3054
rect 2880 -3144 2960 -3106
rect 2880 -3196 2894 -3144
rect 2946 -3196 2960 -3144
rect 2880 -3234 2960 -3196
rect 2880 -3286 2894 -3234
rect 2946 -3286 2960 -3234
rect 2880 -3324 2960 -3286
rect 2880 -3376 2894 -3324
rect 2946 -3376 2960 -3324
rect 2880 -3414 2960 -3376
rect 2880 -3466 2894 -3414
rect 2946 -3466 2960 -3414
rect 2880 -3504 2960 -3466
rect 2880 -3556 2894 -3504
rect 2946 -3556 2960 -3504
rect 2880 -3570 2960 -3556
rect 3260 -3054 3340 -3040
rect 3260 -3106 3274 -3054
rect 3326 -3106 3340 -3054
rect 3260 -3144 3340 -3106
rect 3260 -3196 3274 -3144
rect 3326 -3196 3340 -3144
rect 3260 -3234 3340 -3196
rect 3260 -3286 3274 -3234
rect 3326 -3286 3340 -3234
rect 3260 -3324 3340 -3286
rect 3260 -3376 3274 -3324
rect 3326 -3376 3340 -3324
rect 3260 -3414 3340 -3376
rect 3260 -3466 3274 -3414
rect 3326 -3466 3340 -3414
rect 3260 -3504 3340 -3466
rect 3260 -3556 3274 -3504
rect 3326 -3556 3340 -3504
rect 3260 -3570 3340 -3556
rect 3640 -3054 3720 -3040
rect 3640 -3106 3654 -3054
rect 3706 -3106 3720 -3054
rect 3640 -3144 3720 -3106
rect 3640 -3196 3654 -3144
rect 3706 -3196 3720 -3144
rect 3640 -3234 3720 -3196
rect 3640 -3286 3654 -3234
rect 3706 -3286 3720 -3234
rect 3640 -3324 3720 -3286
rect 3640 -3376 3654 -3324
rect 3706 -3376 3720 -3324
rect 3640 -3414 3720 -3376
rect 3640 -3466 3654 -3414
rect 3706 -3466 3720 -3414
rect 3640 -3504 3720 -3466
rect 3640 -3556 3654 -3504
rect 3706 -3556 3720 -3504
rect 3640 -3570 3720 -3556
rect 4020 -3054 4100 -3040
rect 4020 -3106 4034 -3054
rect 4086 -3106 4100 -3054
rect 4020 -3144 4100 -3106
rect 4020 -3196 4034 -3144
rect 4086 -3196 4100 -3144
rect 4020 -3234 4100 -3196
rect 4020 -3286 4034 -3234
rect 4086 -3286 4100 -3234
rect 4020 -3324 4100 -3286
rect 4020 -3376 4034 -3324
rect 4086 -3376 4100 -3324
rect 4020 -3414 4100 -3376
rect 4020 -3466 4034 -3414
rect 4086 -3466 4100 -3414
rect 4020 -3504 4100 -3466
rect 4020 -3556 4034 -3504
rect 4086 -3556 4100 -3504
rect 4020 -3570 4100 -3556
rect 4130 -4290 4190 -2170
rect 4220 -2290 4480 -2110
rect 4600 -2114 4750 -2110
rect 4600 -2166 4617 -2114
rect 4669 -2166 4681 -2114
rect 4733 -2166 4750 -2114
rect 4600 -2170 4750 -2166
rect 4980 -2114 5130 -2110
rect 4980 -2166 4997 -2114
rect 5049 -2166 5061 -2114
rect 5113 -2166 5130 -2114
rect 4980 -2170 5130 -2166
rect 5360 -2114 5510 -2110
rect 5360 -2166 5377 -2114
rect 5429 -2166 5441 -2114
rect 5493 -2166 5510 -2114
rect 5360 -2170 5510 -2166
rect 5740 -2114 5890 -2110
rect 5740 -2166 5757 -2114
rect 5809 -2166 5821 -2114
rect 5873 -2166 5890 -2114
rect 5740 -2170 5890 -2166
rect 6120 -2114 6470 -2110
rect 6120 -2166 6137 -2114
rect 6189 -2166 6201 -2114
rect 6253 -2166 6470 -2114
rect 6120 -2170 6470 -2166
rect 6500 -2114 6650 -2110
rect 6500 -2166 6517 -2114
rect 6569 -2166 6581 -2114
rect 6633 -2166 6650 -2114
rect 6500 -2170 6650 -2166
rect 6880 -2114 7030 -2110
rect 6880 -2166 6897 -2114
rect 6949 -2166 6961 -2114
rect 7013 -2166 7030 -2114
rect 6880 -2170 7030 -2166
rect 7260 -2114 7410 -2110
rect 7260 -2166 7277 -2114
rect 7329 -2166 7341 -2114
rect 7393 -2166 7410 -2114
rect 7260 -2170 7410 -2166
rect 7640 -2114 7790 -2110
rect 7640 -2166 7657 -2114
rect 7709 -2166 7721 -2114
rect 7773 -2166 7790 -2114
rect 7640 -2170 7790 -2166
rect 8020 -2114 8170 -2110
rect 8020 -2166 8037 -2114
rect 8089 -2166 8101 -2114
rect 8153 -2166 8170 -2114
rect 8020 -2170 8170 -2166
rect 4600 -2234 4750 -2230
rect 4600 -2286 4617 -2234
rect 4669 -2286 4681 -2234
rect 4733 -2286 4750 -2234
rect 4600 -2290 4750 -2286
rect 4980 -2234 5130 -2230
rect 4980 -2286 4997 -2234
rect 5049 -2286 5061 -2234
rect 5113 -2286 5130 -2234
rect 4980 -2290 5130 -2286
rect 5360 -2234 5510 -2230
rect 5360 -2286 5377 -2234
rect 5429 -2286 5441 -2234
rect 5493 -2286 5510 -2234
rect 5360 -2290 5510 -2286
rect 5740 -2234 5890 -2230
rect 5740 -2286 5757 -2234
rect 5809 -2286 5821 -2234
rect 5873 -2286 5890 -2234
rect 5740 -2290 5890 -2286
rect 6120 -2234 6270 -2230
rect 6120 -2286 6137 -2234
rect 6189 -2286 6201 -2234
rect 6253 -2286 6270 -2234
rect 6120 -2290 6270 -2286
rect 4420 -4290 4480 -2290
rect 4780 -3054 4860 -3040
rect 4780 -3106 4794 -3054
rect 4846 -3106 4860 -3054
rect 4780 -3144 4860 -3106
rect 4780 -3196 4794 -3144
rect 4846 -3196 4860 -3144
rect 4780 -3234 4860 -3196
rect 4780 -3286 4794 -3234
rect 4846 -3286 4860 -3234
rect 4780 -3324 4860 -3286
rect 4780 -3376 4794 -3324
rect 4846 -3376 4860 -3324
rect 4780 -3414 4860 -3376
rect 4780 -3466 4794 -3414
rect 4846 -3466 4860 -3414
rect 4780 -3504 4860 -3466
rect 4780 -3556 4794 -3504
rect 4846 -3556 4860 -3504
rect 4780 -3570 4860 -3556
rect 5160 -3054 5240 -3040
rect 5160 -3106 5174 -3054
rect 5226 -3106 5240 -3054
rect 5160 -3144 5240 -3106
rect 5160 -3196 5174 -3144
rect 5226 -3196 5240 -3144
rect 5160 -3234 5240 -3196
rect 5160 -3286 5174 -3234
rect 5226 -3286 5240 -3234
rect 5160 -3324 5240 -3286
rect 5160 -3376 5174 -3324
rect 5226 -3376 5240 -3324
rect 5160 -3414 5240 -3376
rect 5160 -3466 5174 -3414
rect 5226 -3466 5240 -3414
rect 5160 -3504 5240 -3466
rect 5160 -3556 5174 -3504
rect 5226 -3556 5240 -3504
rect 5160 -3570 5240 -3556
rect 5540 -3054 5620 -3040
rect 5540 -3106 5554 -3054
rect 5606 -3106 5620 -3054
rect 5540 -3144 5620 -3106
rect 5540 -3196 5554 -3144
rect 5606 -3196 5620 -3144
rect 5540 -3234 5620 -3196
rect 5540 -3286 5554 -3234
rect 5606 -3286 5620 -3234
rect 5540 -3324 5620 -3286
rect 5540 -3376 5554 -3324
rect 5606 -3376 5620 -3324
rect 5540 -3414 5620 -3376
rect 5540 -3466 5554 -3414
rect 5606 -3466 5620 -3414
rect 5540 -3504 5620 -3466
rect 5540 -3556 5554 -3504
rect 5606 -3556 5620 -3504
rect 5540 -3570 5620 -3556
rect 5920 -3054 6000 -3040
rect 5920 -3106 5934 -3054
rect 5986 -3106 6000 -3054
rect 5920 -3144 6000 -3106
rect 5920 -3196 5934 -3144
rect 5986 -3196 6000 -3144
rect 5920 -3234 6000 -3196
rect 5920 -3286 5934 -3234
rect 5986 -3286 6000 -3234
rect 5920 -3324 6000 -3286
rect 5920 -3376 5934 -3324
rect 5986 -3376 6000 -3324
rect 5920 -3414 6000 -3376
rect 5920 -3466 5934 -3414
rect 5986 -3466 6000 -3414
rect 5920 -3504 6000 -3466
rect 5920 -3556 5934 -3504
rect 5986 -3556 6000 -3504
rect 5920 -3570 6000 -3556
rect 6300 -3054 6380 -3040
rect 6300 -3106 6314 -3054
rect 6366 -3106 6380 -3054
rect 6300 -3144 6380 -3106
rect 6300 -3196 6314 -3144
rect 6366 -3196 6380 -3144
rect 6300 -3234 6380 -3196
rect 6300 -3286 6314 -3234
rect 6366 -3286 6380 -3234
rect 6300 -3324 6380 -3286
rect 6300 -3376 6314 -3324
rect 6366 -3376 6380 -3324
rect 6300 -3414 6380 -3376
rect 6300 -3466 6314 -3414
rect 6366 -3466 6380 -3414
rect 6300 -3504 6380 -3466
rect 6300 -3556 6314 -3504
rect 6366 -3556 6380 -3504
rect 6300 -3570 6380 -3556
rect 6410 -4290 6470 -2170
rect 6500 -2234 6650 -2230
rect 6500 -2286 6517 -2234
rect 6569 -2286 6581 -2234
rect 6633 -2286 6650 -2234
rect 6500 -2290 6650 -2286
rect 6880 -2234 7030 -2230
rect 6880 -2286 6897 -2234
rect 6949 -2286 6961 -2234
rect 7013 -2286 7030 -2234
rect 6880 -2290 7030 -2286
rect 7260 -2234 7410 -2230
rect 7260 -2286 7277 -2234
rect 7329 -2286 7341 -2234
rect 7393 -2286 7410 -2234
rect 7260 -2290 7410 -2286
rect 7640 -2234 7790 -2230
rect 7640 -2286 7657 -2234
rect 7709 -2286 7721 -2234
rect 7773 -2286 7790 -2234
rect 7640 -2290 7790 -2286
rect 8020 -2234 8170 -2230
rect 8020 -2286 8037 -2234
rect 8089 -2286 8101 -2234
rect 8153 -2286 8170 -2234
rect 8020 -2290 8170 -2286
rect 8370 -2290 8660 -2110
rect 6680 -3054 6760 -3040
rect 6680 -3106 6694 -3054
rect 6746 -3106 6760 -3054
rect 6680 -3144 6760 -3106
rect 6680 -3196 6694 -3144
rect 6746 -3196 6760 -3144
rect 6680 -3234 6760 -3196
rect 6680 -3286 6694 -3234
rect 6746 -3286 6760 -3234
rect 6680 -3324 6760 -3286
rect 6680 -3376 6694 -3324
rect 6746 -3376 6760 -3324
rect 6680 -3414 6760 -3376
rect 6680 -3466 6694 -3414
rect 6746 -3466 6760 -3414
rect 6680 -3504 6760 -3466
rect 6680 -3556 6694 -3504
rect 6746 -3556 6760 -3504
rect 6680 -3570 6760 -3556
rect 7060 -3054 7140 -3040
rect 7060 -3106 7074 -3054
rect 7126 -3106 7140 -3054
rect 7060 -3144 7140 -3106
rect 7060 -3196 7074 -3144
rect 7126 -3196 7140 -3144
rect 7060 -3234 7140 -3196
rect 7060 -3286 7074 -3234
rect 7126 -3286 7140 -3234
rect 7060 -3324 7140 -3286
rect 7060 -3376 7074 -3324
rect 7126 -3376 7140 -3324
rect 7060 -3414 7140 -3376
rect 7060 -3466 7074 -3414
rect 7126 -3466 7140 -3414
rect 7060 -3504 7140 -3466
rect 7060 -3556 7074 -3504
rect 7126 -3556 7140 -3504
rect 7060 -3570 7140 -3556
rect 7440 -3054 7520 -3040
rect 7440 -3106 7454 -3054
rect 7506 -3106 7520 -3054
rect 7440 -3144 7520 -3106
rect 7440 -3196 7454 -3144
rect 7506 -3196 7520 -3144
rect 7440 -3234 7520 -3196
rect 7440 -3286 7454 -3234
rect 7506 -3286 7520 -3234
rect 7440 -3324 7520 -3286
rect 7440 -3376 7454 -3324
rect 7506 -3376 7520 -3324
rect 7440 -3414 7520 -3376
rect 7440 -3466 7454 -3414
rect 7506 -3466 7520 -3414
rect 7440 -3504 7520 -3466
rect 7440 -3556 7454 -3504
rect 7506 -3556 7520 -3504
rect 7440 -3570 7520 -3556
rect 7820 -3054 7900 -3040
rect 7820 -3106 7834 -3054
rect 7886 -3106 7900 -3054
rect 7820 -3144 7900 -3106
rect 7820 -3196 7834 -3144
rect 7886 -3196 7900 -3144
rect 7820 -3234 7900 -3196
rect 7820 -3286 7834 -3234
rect 7886 -3286 7900 -3234
rect 7820 -3324 7900 -3286
rect 7820 -3376 7834 -3324
rect 7886 -3376 7900 -3324
rect 7820 -3414 7900 -3376
rect 7820 -3466 7834 -3414
rect 7886 -3466 7900 -3414
rect 7820 -3504 7900 -3466
rect 7820 -3556 7834 -3504
rect 7886 -3556 7900 -3504
rect 7820 -3570 7900 -3556
rect 8200 -3054 8280 -3040
rect 8200 -3106 8214 -3054
rect 8266 -3106 8280 -3054
rect 8200 -3144 8280 -3106
rect 8200 -3196 8214 -3144
rect 8266 -3196 8280 -3144
rect 8200 -3234 8280 -3196
rect 8200 -3286 8214 -3234
rect 8266 -3286 8280 -3234
rect 8200 -3324 8280 -3286
rect 8200 -3376 8214 -3324
rect 8266 -3376 8280 -3324
rect 8200 -3414 8280 -3376
rect 8200 -3466 8214 -3414
rect 8266 -3466 8280 -3414
rect 8200 -3504 8280 -3466
rect 8200 -3556 8214 -3504
rect 8266 -3556 8280 -3504
rect 8200 -3570 8280 -3556
rect 8600 -4290 8660 -2290
rect -250 -4346 -236 -4294
rect -184 -4346 -170 -4294
rect -250 -4684 -170 -4346
rect -250 -4736 -236 -4684
rect -184 -4736 -170 -4684
rect -250 -4764 -170 -4736
rect -250 -4816 -236 -4764
rect -184 -4816 -170 -4764
rect -250 -4820 -170 -4816
rect 10 -4410 300 -4290
rect 420 -4294 570 -4290
rect 420 -4346 437 -4294
rect 489 -4346 501 -4294
rect 553 -4346 570 -4294
rect 420 -4350 570 -4346
rect 800 -4294 950 -4290
rect 800 -4346 817 -4294
rect 869 -4346 881 -4294
rect 933 -4346 950 -4294
rect 800 -4350 950 -4346
rect 1180 -4294 1330 -4290
rect 1180 -4346 1197 -4294
rect 1249 -4346 1261 -4294
rect 1313 -4346 1330 -4294
rect 1180 -4350 1330 -4346
rect 1560 -4294 1710 -4290
rect 1560 -4346 1577 -4294
rect 1629 -4346 1641 -4294
rect 1693 -4346 1710 -4294
rect 1560 -4350 1710 -4346
rect 1940 -4294 2090 -4290
rect 1940 -4346 1957 -4294
rect 2009 -4346 2021 -4294
rect 2073 -4346 2090 -4294
rect 1940 -4350 2090 -4346
rect 2320 -4294 2470 -4290
rect 2320 -4346 2337 -4294
rect 2389 -4346 2401 -4294
rect 2453 -4346 2470 -4294
rect 2320 -4350 2470 -4346
rect 2700 -4294 2850 -4290
rect 2700 -4346 2717 -4294
rect 2769 -4346 2781 -4294
rect 2833 -4346 2850 -4294
rect 2700 -4350 2850 -4346
rect 3080 -4294 3230 -4290
rect 3080 -4346 3097 -4294
rect 3149 -4346 3161 -4294
rect 3213 -4346 3230 -4294
rect 3080 -4350 3230 -4346
rect 3460 -4294 3610 -4290
rect 3460 -4346 3477 -4294
rect 3529 -4346 3541 -4294
rect 3593 -4346 3610 -4294
rect 3460 -4350 3610 -4346
rect 3840 -4294 4190 -4290
rect 3840 -4346 3857 -4294
rect 3909 -4346 3921 -4294
rect 3973 -4346 4024 -4294
rect 4076 -4346 4124 -4294
rect 4176 -4346 4190 -4294
rect 3840 -4350 4190 -4346
rect 4220 -4410 4480 -4290
rect 4600 -4294 4750 -4290
rect 4600 -4346 4617 -4294
rect 4669 -4346 4681 -4294
rect 4733 -4346 4750 -4294
rect 4600 -4350 4750 -4346
rect 4980 -4294 5130 -4290
rect 4980 -4346 4997 -4294
rect 5049 -4346 5061 -4294
rect 5113 -4346 5130 -4294
rect 4980 -4350 5130 -4346
rect 5360 -4294 5510 -4290
rect 5360 -4346 5377 -4294
rect 5429 -4346 5441 -4294
rect 5493 -4346 5510 -4294
rect 5360 -4350 5510 -4346
rect 5740 -4294 5890 -4290
rect 5740 -4346 5757 -4294
rect 5809 -4346 5821 -4294
rect 5873 -4346 5890 -4294
rect 5740 -4350 5890 -4346
rect 6120 -4294 6470 -4290
rect 6120 -4346 6137 -4294
rect 6189 -4346 6201 -4294
rect 6253 -4346 6314 -4294
rect 6366 -4346 6404 -4294
rect 6456 -4346 6470 -4294
rect 6120 -4350 6470 -4346
rect 6500 -4294 6650 -4290
rect 6500 -4346 6517 -4294
rect 6569 -4346 6581 -4294
rect 6633 -4346 6650 -4294
rect 6500 -4350 6650 -4346
rect 6880 -4294 7030 -4290
rect 6880 -4346 6897 -4294
rect 6949 -4346 6961 -4294
rect 7013 -4346 7030 -4294
rect 6880 -4350 7030 -4346
rect 7260 -4294 7410 -4290
rect 7260 -4346 7277 -4294
rect 7329 -4346 7341 -4294
rect 7393 -4346 7410 -4294
rect 7260 -4350 7410 -4346
rect 7640 -4294 7790 -4290
rect 7640 -4346 7657 -4294
rect 7709 -4346 7721 -4294
rect 7773 -4346 7790 -4294
rect 7640 -4350 7790 -4346
rect 8020 -4294 8170 -4290
rect 8020 -4346 8037 -4294
rect 8089 -4346 8101 -4294
rect 8153 -4346 8170 -4294
rect 8020 -4350 8170 -4346
rect 8380 -4410 8660 -4290
rect 10 -4730 8660 -4410
rect 8690 -2034 8770 -2030
rect 8690 -2086 8704 -2034
rect 8756 -2086 8770 -2034
rect 8690 -2114 8770 -2086
rect 8690 -2166 8704 -2114
rect 8756 -2166 8770 -2114
rect 8690 -4294 8770 -2166
rect 8690 -4346 8704 -4294
rect 8756 -4346 8770 -4294
rect 8690 -4374 8770 -4346
rect 8690 -4426 8704 -4374
rect 8756 -4426 8770 -4374
rect 10 -5320 370 -4730
rect 2130 -5320 2490 -4730
rect 5860 -5320 6220 -4730
rect 8220 -5320 8580 -4730
rect 8690 -5004 8770 -4426
rect 8690 -5056 8704 -5004
rect 8756 -5056 8770 -5004
rect 8690 -5084 8770 -5056
rect 8690 -5136 8704 -5084
rect 8756 -5136 8770 -5084
rect 8690 -5150 8770 -5136
<< via1 >>
rect 8764 5034 8816 5086
rect 8844 5034 8896 5086
rect 2144 4714 2196 4766
rect 2224 4714 2276 4766
rect 1934 4374 1986 4426
rect 2014 4374 2066 4426
rect 437 4254 489 4306
rect 501 4254 553 4306
rect 817 4254 869 4306
rect 881 4254 933 4306
rect 1197 4254 1249 4306
rect 1261 4254 1313 4306
rect 1577 4254 1629 4306
rect 1641 4254 1693 4306
rect 1957 4254 2009 4306
rect 2021 4254 2073 4306
rect -96 2274 -44 2326
rect 614 3474 666 3526
rect 614 3384 666 3436
rect 614 3294 666 3346
rect 614 3204 666 3256
rect 614 3114 666 3166
rect 614 3024 666 3076
rect 994 3474 1046 3526
rect 994 3384 1046 3436
rect 994 3294 1046 3346
rect 994 3204 1046 3256
rect 994 3114 1046 3166
rect 994 3024 1046 3076
rect 1374 3474 1426 3526
rect 1374 3384 1426 3436
rect 1374 3294 1426 3346
rect 1374 3204 1426 3256
rect 1374 3114 1426 3166
rect 1374 3024 1426 3076
rect 1754 3474 1806 3526
rect 1754 3384 1806 3436
rect 1754 3294 1806 3346
rect 1754 3204 1806 3256
rect 1754 3114 1806 3166
rect 1754 3024 1806 3076
rect 2134 3474 2186 3526
rect 2134 3384 2186 3436
rect 2134 3294 2186 3346
rect 2134 3204 2186 3256
rect 2134 3114 2186 3166
rect 2134 3024 2186 3076
rect 2334 4374 2386 4426
rect 2434 4374 2486 4426
rect 2337 4254 2389 4306
rect 2401 4254 2453 4306
rect 2717 4254 2769 4306
rect 2781 4254 2833 4306
rect 3097 4254 3149 4306
rect 3161 4254 3213 4306
rect 3477 4254 3529 4306
rect 3541 4254 3593 4306
rect 3857 4254 3909 4306
rect 3921 4254 3973 4306
rect 2514 3474 2566 3526
rect 2514 3384 2566 3436
rect 2514 3294 2566 3346
rect 2514 3204 2566 3256
rect 2514 3114 2566 3166
rect 2514 3024 2566 3076
rect 2894 3474 2946 3526
rect 2894 3384 2946 3436
rect 2894 3294 2946 3346
rect 2894 3204 2946 3256
rect 2894 3114 2946 3166
rect 2894 3024 2946 3076
rect 3274 3474 3326 3526
rect 3274 3384 3326 3436
rect 3274 3294 3326 3346
rect 3274 3204 3326 3256
rect 3274 3114 3326 3166
rect 3274 3024 3326 3076
rect 3654 3474 3706 3526
rect 3654 3384 3706 3436
rect 3654 3294 3706 3346
rect 3654 3204 3706 3256
rect 3654 3114 3706 3166
rect 3654 3024 3706 3076
rect 4034 3474 4086 3526
rect 4034 3384 4086 3436
rect 4034 3294 4086 3346
rect 4034 3204 4086 3256
rect 4034 3114 4086 3166
rect 4034 3024 4086 3076
rect -96 2194 -44 2246
rect 437 2194 489 2246
rect 501 2194 553 2246
rect 817 2194 869 2246
rect 881 2194 933 2246
rect 1197 2194 1249 2246
rect 1261 2194 1313 2246
rect 1577 2194 1629 2246
rect 1641 2194 1693 2246
rect 1957 2194 2009 2246
rect 2021 2194 2073 2246
rect 2337 2194 2389 2246
rect 2401 2194 2453 2246
rect 2717 2194 2769 2246
rect 2781 2194 2833 2246
rect 3097 2194 3149 2246
rect 3161 2194 3213 2246
rect 3477 2194 3529 2246
rect 3541 2194 3593 2246
rect 3857 2194 3909 2246
rect 3921 2194 3973 2246
rect 4524 4264 4576 4316
rect 4614 4259 4666 4311
rect 4685 4254 4737 4306
rect 4997 4254 5049 4306
rect 5061 4254 5113 4306
rect 5377 4254 5429 4306
rect 5441 4254 5493 4306
rect 5757 4254 5809 4306
rect 5821 4254 5873 4306
rect 6137 4254 6189 4306
rect 6201 4254 6253 4306
rect 6517 4254 6569 4306
rect 6581 4254 6633 4306
rect 6897 4254 6949 4306
rect 6961 4254 7013 4306
rect 7277 4254 7329 4306
rect 7341 4254 7393 4306
rect 7657 4254 7709 4306
rect 7721 4254 7773 4306
rect 8037 4254 8089 4306
rect 8101 4254 8153 4306
rect 437 2074 489 2126
rect 501 2074 553 2126
rect 817 2074 869 2126
rect 881 2074 933 2126
rect 1197 2074 1249 2126
rect 1261 2074 1313 2126
rect 1577 2074 1629 2126
rect 1641 2074 1693 2126
rect 1957 2074 2009 2126
rect 2021 2074 2073 2126
rect -96 1744 -44 1796
rect -96 1654 -44 1706
rect 614 1324 666 1376
rect 614 1234 666 1286
rect 614 1144 666 1196
rect 614 1054 666 1106
rect 614 964 666 1016
rect 614 874 666 926
rect 994 1324 1046 1376
rect 994 1234 1046 1286
rect 994 1144 1046 1196
rect 994 1054 1046 1106
rect 994 964 1046 1016
rect 994 874 1046 926
rect 1374 1324 1426 1376
rect 1374 1234 1426 1286
rect 1374 1144 1426 1196
rect 1374 1054 1426 1106
rect 1374 964 1426 1016
rect 1374 874 1426 926
rect 1754 1324 1806 1376
rect 1754 1234 1806 1286
rect 1754 1144 1806 1196
rect 1754 1054 1806 1106
rect 1754 964 1806 1016
rect 1754 874 1806 926
rect 2134 1324 2186 1376
rect 2134 1234 2186 1286
rect 2134 1144 2186 1196
rect 2134 1054 2186 1106
rect 2134 964 2186 1016
rect 2134 874 2186 926
rect 2337 2074 2389 2126
rect 2401 2074 2453 2126
rect 2717 2074 2769 2126
rect 2781 2074 2833 2126
rect 3097 2074 3149 2126
rect 3161 2074 3213 2126
rect 3477 2074 3529 2126
rect 3541 2074 3593 2126
rect 3857 2074 3909 2126
rect 3921 2074 3973 2126
rect 2514 1324 2566 1376
rect 2514 1234 2566 1286
rect 2514 1144 2566 1196
rect 2514 1054 2566 1106
rect 2514 964 2566 1016
rect 2514 874 2566 926
rect 2894 1324 2946 1376
rect 2894 1234 2946 1286
rect 2894 1144 2946 1196
rect 2894 1054 2946 1106
rect 2894 964 2946 1016
rect 2894 874 2946 926
rect 3274 1324 3326 1376
rect 3274 1234 3326 1286
rect 3274 1144 3326 1196
rect 3274 1054 3326 1106
rect 3274 964 3326 1016
rect 3274 874 3326 926
rect 3654 1324 3706 1376
rect 3654 1234 3706 1286
rect 3654 1144 3706 1196
rect 3654 1054 3706 1106
rect 3654 964 3706 1016
rect 3654 874 3706 926
rect 4034 1324 4086 1376
rect 4034 1234 4086 1286
rect 4034 1144 4086 1196
rect 4034 1054 4086 1106
rect 4034 964 4086 1016
rect 4034 874 4086 926
rect 4234 2084 4286 2136
rect 4324 2084 4376 2136
rect 4794 3474 4846 3526
rect 4794 3384 4846 3436
rect 4794 3294 4846 3346
rect 4794 3204 4846 3256
rect 4794 3114 4846 3166
rect 4794 3024 4846 3076
rect 5174 3474 5226 3526
rect 5174 3384 5226 3436
rect 5174 3294 5226 3346
rect 5174 3204 5226 3256
rect 5174 3114 5226 3166
rect 5174 3024 5226 3076
rect 5554 3474 5606 3526
rect 5554 3384 5606 3436
rect 5554 3294 5606 3346
rect 5554 3204 5606 3256
rect 5554 3114 5606 3166
rect 5554 3024 5606 3076
rect 5934 3474 5986 3526
rect 5934 3384 5986 3436
rect 5934 3294 5986 3346
rect 5934 3204 5986 3256
rect 5934 3114 5986 3166
rect 5934 3024 5986 3076
rect 6314 3474 6366 3526
rect 6314 3384 6366 3436
rect 6314 3294 6366 3346
rect 6314 3204 6366 3256
rect 6314 3114 6366 3166
rect 6314 3024 6366 3076
rect 6694 3474 6746 3526
rect 6694 3384 6746 3436
rect 6694 3294 6746 3346
rect 6694 3204 6746 3256
rect 6694 3114 6746 3166
rect 6694 3024 6746 3076
rect 7074 3474 7126 3526
rect 7074 3384 7126 3436
rect 7074 3294 7126 3346
rect 7074 3204 7126 3256
rect 7074 3114 7126 3166
rect 7074 3024 7126 3076
rect 7454 3474 7506 3526
rect 7454 3384 7506 3436
rect 7454 3294 7506 3346
rect 7454 3204 7506 3256
rect 7454 3114 7506 3166
rect 7454 3024 7506 3076
rect 7834 3474 7886 3526
rect 7834 3384 7886 3436
rect 7834 3294 7886 3346
rect 7834 3204 7886 3256
rect 7834 3114 7886 3166
rect 7834 3024 7886 3076
rect 8214 3474 8266 3526
rect 8214 3384 8266 3436
rect 8214 3294 8266 3346
rect 8214 3204 8266 3256
rect 8214 3114 8266 3166
rect 8214 3024 8266 3076
rect 4617 2194 4669 2246
rect 4681 2194 4733 2246
rect 4997 2194 5049 2246
rect 5061 2194 5113 2246
rect 5377 2194 5429 2246
rect 5441 2194 5493 2246
rect 5757 2194 5809 2246
rect 5821 2194 5873 2246
rect 6137 2194 6189 2246
rect 6201 2194 6253 2246
rect 6517 2194 6569 2246
rect 6581 2194 6633 2246
rect 6897 2194 6949 2246
rect 6961 2194 7013 2246
rect 7277 2194 7329 2246
rect 7341 2194 7393 2246
rect 7657 2194 7709 2246
rect 7721 2194 7773 2246
rect 8037 2194 8089 2246
rect 8101 2194 8153 2246
rect 4617 2074 4669 2126
rect 4681 2074 4733 2126
rect 4997 2074 5049 2126
rect 5061 2074 5113 2126
rect 5377 2074 5429 2126
rect 5441 2074 5493 2126
rect 5757 2074 5809 2126
rect 5821 2074 5873 2126
rect 6137 2074 6189 2126
rect 6201 2074 6253 2126
rect 6517 2074 6569 2126
rect 6581 2074 6633 2126
rect 6897 2074 6949 2126
rect 6961 2074 7013 2126
rect 7277 2074 7329 2126
rect 7341 2074 7393 2126
rect 7657 2074 7709 2126
rect 7721 2074 7773 2126
rect 8037 2074 8089 2126
rect 8101 2074 8153 2126
rect 437 14 489 66
rect 501 14 553 66
rect 817 14 869 66
rect 881 14 933 66
rect 1197 14 1249 66
rect 1261 14 1313 66
rect 1577 14 1629 66
rect 1641 14 1693 66
rect 1957 14 2009 66
rect 2021 14 2073 66
rect 2337 14 2389 66
rect 2401 14 2453 66
rect 2717 14 2769 66
rect 2781 14 2833 66
rect 3097 14 3149 66
rect 3161 14 3213 66
rect 3477 14 3529 66
rect 3541 14 3593 66
rect 3857 14 3909 66
rect 3921 14 3973 66
rect 4794 1324 4846 1376
rect 4794 1234 4846 1286
rect 4794 1144 4846 1196
rect 4794 1054 4846 1106
rect 4794 964 4846 1016
rect 4794 874 4846 926
rect 5174 1324 5226 1376
rect 5174 1234 5226 1286
rect 5174 1144 5226 1196
rect 5174 1054 5226 1106
rect 5174 964 5226 1016
rect 5174 874 5226 926
rect 5554 1324 5606 1376
rect 5554 1234 5606 1286
rect 5554 1144 5606 1196
rect 5554 1054 5606 1106
rect 5554 964 5606 1016
rect 5554 874 5606 926
rect 5934 1324 5986 1376
rect 5934 1234 5986 1286
rect 5934 1144 5986 1196
rect 5934 1054 5986 1106
rect 5934 964 5986 1016
rect 5934 874 5986 926
rect 6314 1324 6366 1376
rect 6314 1234 6366 1286
rect 6314 1144 6366 1196
rect 6314 1054 6366 1106
rect 6314 964 6366 1016
rect 6314 874 6366 926
rect 6694 1324 6746 1376
rect 6694 1234 6746 1286
rect 6694 1144 6746 1196
rect 6694 1054 6746 1106
rect 6694 964 6746 1016
rect 6694 874 6746 926
rect 7074 1324 7126 1376
rect 7074 1234 7126 1286
rect 7074 1144 7126 1196
rect 7074 1054 7126 1106
rect 7074 964 7126 1016
rect 7074 874 7126 926
rect 7454 1324 7506 1376
rect 7454 1234 7506 1286
rect 7454 1144 7506 1196
rect 7454 1054 7506 1106
rect 7454 964 7506 1016
rect 7454 874 7506 926
rect 7834 1324 7886 1376
rect 7834 1234 7886 1286
rect 7834 1144 7886 1196
rect 7834 1054 7886 1106
rect 7834 964 7886 1016
rect 7834 874 7886 926
rect 8214 1324 8266 1376
rect 8214 1234 8266 1286
rect 8214 1144 8266 1196
rect 8214 1054 8266 1106
rect 8214 964 8266 1016
rect 8214 874 8266 926
rect 8844 4254 8896 4306
rect 8844 4174 8896 4226
rect 8844 2074 8896 2126
rect 8844 1994 8896 2046
rect 4617 14 4669 66
rect 4681 14 4733 66
rect 4997 14 5049 66
rect 5061 14 5113 66
rect 5377 14 5429 66
rect 5441 14 5493 66
rect 5757 14 5809 66
rect 5821 14 5873 66
rect 6137 14 6189 66
rect 6201 14 6253 66
rect 6517 14 6569 66
rect 6581 14 6633 66
rect 6897 14 6949 66
rect 6961 14 7013 66
rect 7277 14 7329 66
rect 7341 14 7393 66
rect 7657 14 7709 66
rect 7721 14 7773 66
rect 8037 14 8089 66
rect 8101 14 8153 66
rect 437 -106 489 -54
rect 501 -106 553 -54
rect 817 -106 869 -54
rect 881 -106 933 -54
rect 1197 -106 1249 -54
rect 1261 -106 1313 -54
rect 1577 -106 1629 -54
rect 1641 -106 1693 -54
rect 1957 -106 2009 -54
rect 2021 -106 2073 -54
rect 2337 -106 2389 -54
rect 2401 -106 2453 -54
rect 2717 -106 2769 -54
rect 2781 -106 2833 -54
rect 3097 -106 3149 -54
rect 3161 -106 3213 -54
rect 3477 -106 3529 -54
rect 3541 -106 3593 -54
rect 3857 -106 3909 -54
rect 3921 -106 3973 -54
rect 4617 -106 4669 -54
rect 4681 -106 4733 -54
rect 4997 -106 5049 -54
rect 5061 -106 5113 -54
rect 5377 -106 5429 -54
rect 5441 -106 5493 -54
rect 5757 -106 5809 -54
rect 5821 -106 5873 -54
rect 6137 -106 6189 -54
rect 6201 -106 6253 -54
rect 6517 -106 6569 -54
rect 6581 -106 6633 -54
rect 6897 -106 6949 -54
rect 6961 -106 7013 -54
rect 7277 -106 7329 -54
rect 7341 -106 7393 -54
rect 7657 -106 7709 -54
rect 7721 -106 7773 -54
rect 8037 -106 8089 -54
rect 8101 -106 8153 -54
rect -236 -2086 -184 -2034
rect 614 -916 666 -864
rect 614 -1006 666 -954
rect 614 -1096 666 -1044
rect 614 -1186 666 -1134
rect 614 -1276 666 -1224
rect 614 -1366 666 -1314
rect 994 -916 1046 -864
rect 994 -1006 1046 -954
rect 994 -1096 1046 -1044
rect 994 -1186 1046 -1134
rect 994 -1276 1046 -1224
rect 994 -1366 1046 -1314
rect 1374 -916 1426 -864
rect 1374 -1006 1426 -954
rect 1374 -1096 1426 -1044
rect 1374 -1186 1426 -1134
rect 1374 -1276 1426 -1224
rect 1374 -1366 1426 -1314
rect 1754 -916 1806 -864
rect 1754 -1006 1806 -954
rect 1754 -1096 1806 -1044
rect 1754 -1186 1806 -1134
rect 1754 -1276 1806 -1224
rect 1754 -1366 1806 -1314
rect 2134 -916 2186 -864
rect 2134 -1006 2186 -954
rect 2134 -1096 2186 -1044
rect 2134 -1186 2186 -1134
rect 2134 -1276 2186 -1224
rect 2134 -1366 2186 -1314
rect 2514 -916 2566 -864
rect 2514 -1006 2566 -954
rect 2514 -1096 2566 -1044
rect 2514 -1186 2566 -1134
rect 2514 -1276 2566 -1224
rect 2514 -1366 2566 -1314
rect 2894 -916 2946 -864
rect 2894 -1006 2946 -954
rect 2894 -1096 2946 -1044
rect 2894 -1186 2946 -1134
rect 2894 -1276 2946 -1224
rect 2894 -1366 2946 -1314
rect 3274 -916 3326 -864
rect 3274 -1006 3326 -954
rect 3274 -1096 3326 -1044
rect 3274 -1186 3326 -1134
rect 3274 -1276 3326 -1224
rect 3274 -1366 3326 -1314
rect 3654 -916 3706 -864
rect 3654 -1006 3706 -954
rect 3654 -1096 3706 -1044
rect 3654 -1186 3706 -1134
rect 3654 -1276 3706 -1224
rect 3654 -1366 3706 -1314
rect 4034 -916 4086 -864
rect 4034 -1006 4086 -954
rect 4034 -1096 4086 -1044
rect 4034 -1186 4086 -1134
rect 4034 -1276 4086 -1224
rect 4034 -1366 4086 -1314
rect 4794 -916 4846 -864
rect 4794 -1006 4846 -954
rect 4794 -1096 4846 -1044
rect 4794 -1186 4846 -1134
rect 4794 -1276 4846 -1224
rect 4794 -1366 4846 -1314
rect 5174 -916 5226 -864
rect 5174 -1006 5226 -954
rect 5174 -1096 5226 -1044
rect 5174 -1186 5226 -1134
rect 5174 -1276 5226 -1224
rect 5174 -1366 5226 -1314
rect 5554 -916 5606 -864
rect 5554 -1006 5606 -954
rect 5554 -1096 5606 -1044
rect 5554 -1186 5606 -1134
rect 5554 -1276 5606 -1224
rect 5554 -1366 5606 -1314
rect 5934 -916 5986 -864
rect 5934 -1006 5986 -954
rect 5934 -1096 5986 -1044
rect 5934 -1186 5986 -1134
rect 5934 -1276 5986 -1224
rect 5934 -1366 5986 -1314
rect 6314 -916 6366 -864
rect 6314 -1006 6366 -954
rect 6314 -1096 6366 -1044
rect 6314 -1186 6366 -1134
rect 6314 -1276 6366 -1224
rect 6314 -1366 6366 -1314
rect 6694 -916 6746 -864
rect 6694 -1006 6746 -954
rect 6694 -1096 6746 -1044
rect 6694 -1186 6746 -1134
rect 6694 -1276 6746 -1224
rect 6694 -1366 6746 -1314
rect 7074 -916 7126 -864
rect 7074 -1006 7126 -954
rect 7074 -1096 7126 -1044
rect 7074 -1186 7126 -1134
rect 7074 -1276 7126 -1224
rect 7074 -1366 7126 -1314
rect 7454 -916 7506 -864
rect 7454 -1006 7506 -954
rect 7454 -1096 7506 -1044
rect 7454 -1186 7506 -1134
rect 7454 -1276 7506 -1224
rect 7454 -1366 7506 -1314
rect 7834 -916 7886 -864
rect 7834 -1006 7886 -954
rect 7834 -1096 7886 -1044
rect 7834 -1186 7886 -1134
rect 7834 -1276 7886 -1224
rect 7834 -1366 7886 -1314
rect 8214 -916 8266 -864
rect 8214 -1006 8266 -954
rect 8214 -1096 8266 -1044
rect 8214 -1186 8266 -1134
rect 8214 -1276 8266 -1224
rect 8214 -1366 8266 -1314
rect -236 -2166 -184 -2114
rect 437 -2166 489 -2114
rect 501 -2166 553 -2114
rect 817 -2166 869 -2114
rect 881 -2166 933 -2114
rect 1197 -2166 1249 -2114
rect 1261 -2166 1313 -2114
rect 1577 -2166 1629 -2114
rect 1641 -2166 1693 -2114
rect 1957 -2166 2009 -2114
rect 2021 -2166 2073 -2114
rect 2337 -2166 2389 -2114
rect 2401 -2166 2453 -2114
rect 2717 -2166 2769 -2114
rect 2781 -2166 2833 -2114
rect 3097 -2166 3149 -2114
rect 3161 -2166 3213 -2114
rect 3477 -2166 3529 -2114
rect 3541 -2166 3593 -2114
rect 3857 -2166 3909 -2114
rect 3921 -2166 3973 -2114
rect 4004 -2166 4056 -2114
rect 437 -2286 489 -2234
rect 501 -2286 553 -2234
rect 817 -2286 869 -2234
rect 881 -2286 933 -2234
rect 1197 -2286 1249 -2234
rect 1261 -2286 1313 -2234
rect 1577 -2286 1629 -2234
rect 1641 -2286 1693 -2234
rect 1957 -2286 2009 -2234
rect 2021 -2286 2073 -2234
rect 2337 -2286 2389 -2234
rect 2401 -2286 2453 -2234
rect 2717 -2286 2769 -2234
rect 2781 -2286 2833 -2234
rect 3097 -2286 3149 -2234
rect 3161 -2286 3213 -2234
rect 3477 -2286 3529 -2234
rect 3541 -2286 3593 -2234
rect 3857 -2286 3909 -2234
rect 3921 -2286 3973 -2234
rect -236 -4266 -184 -4214
rect 614 -3106 666 -3054
rect 614 -3196 666 -3144
rect 614 -3286 666 -3234
rect 614 -3376 666 -3324
rect 614 -3466 666 -3414
rect 614 -3556 666 -3504
rect 994 -3106 1046 -3054
rect 994 -3196 1046 -3144
rect 994 -3286 1046 -3234
rect 994 -3376 1046 -3324
rect 994 -3466 1046 -3414
rect 994 -3556 1046 -3504
rect 1374 -3106 1426 -3054
rect 1374 -3196 1426 -3144
rect 1374 -3286 1426 -3234
rect 1374 -3376 1426 -3324
rect 1374 -3466 1426 -3414
rect 1374 -3556 1426 -3504
rect 1754 -3106 1806 -3054
rect 1754 -3196 1806 -3144
rect 1754 -3286 1806 -3234
rect 1754 -3376 1806 -3324
rect 1754 -3466 1806 -3414
rect 1754 -3556 1806 -3504
rect 2134 -3106 2186 -3054
rect 2134 -3196 2186 -3144
rect 2134 -3286 2186 -3234
rect 2134 -3376 2186 -3324
rect 2134 -3466 2186 -3414
rect 2134 -3556 2186 -3504
rect 2514 -3106 2566 -3054
rect 2514 -3196 2566 -3144
rect 2514 -3286 2566 -3234
rect 2514 -3376 2566 -3324
rect 2514 -3466 2566 -3414
rect 2514 -3556 2566 -3504
rect 2894 -3106 2946 -3054
rect 2894 -3196 2946 -3144
rect 2894 -3286 2946 -3234
rect 2894 -3376 2946 -3324
rect 2894 -3466 2946 -3414
rect 2894 -3556 2946 -3504
rect 3274 -3106 3326 -3054
rect 3274 -3196 3326 -3144
rect 3274 -3286 3326 -3234
rect 3274 -3376 3326 -3324
rect 3274 -3466 3326 -3414
rect 3274 -3556 3326 -3504
rect 3654 -3106 3706 -3054
rect 3654 -3196 3706 -3144
rect 3654 -3286 3706 -3234
rect 3654 -3376 3706 -3324
rect 3654 -3466 3706 -3414
rect 3654 -3556 3706 -3504
rect 4034 -3106 4086 -3054
rect 4034 -3196 4086 -3144
rect 4034 -3286 4086 -3234
rect 4034 -3376 4086 -3324
rect 4034 -3466 4086 -3414
rect 4034 -3556 4086 -3504
rect 4617 -2166 4669 -2114
rect 4681 -2166 4733 -2114
rect 4997 -2166 5049 -2114
rect 5061 -2166 5113 -2114
rect 5377 -2166 5429 -2114
rect 5441 -2166 5493 -2114
rect 5757 -2166 5809 -2114
rect 5821 -2166 5873 -2114
rect 6137 -2166 6189 -2114
rect 6201 -2166 6253 -2114
rect 6517 -2166 6569 -2114
rect 6581 -2166 6633 -2114
rect 6897 -2166 6949 -2114
rect 6961 -2166 7013 -2114
rect 7277 -2166 7329 -2114
rect 7341 -2166 7393 -2114
rect 7657 -2166 7709 -2114
rect 7721 -2166 7773 -2114
rect 8037 -2166 8089 -2114
rect 8101 -2166 8153 -2114
rect 4617 -2286 4669 -2234
rect 4681 -2286 4733 -2234
rect 4997 -2286 5049 -2234
rect 5061 -2286 5113 -2234
rect 5377 -2286 5429 -2234
rect 5441 -2286 5493 -2234
rect 5757 -2286 5809 -2234
rect 5821 -2286 5873 -2234
rect 6137 -2286 6189 -2234
rect 6201 -2286 6253 -2234
rect 4794 -3106 4846 -3054
rect 4794 -3196 4846 -3144
rect 4794 -3286 4846 -3234
rect 4794 -3376 4846 -3324
rect 4794 -3466 4846 -3414
rect 4794 -3556 4846 -3504
rect 5174 -3106 5226 -3054
rect 5174 -3196 5226 -3144
rect 5174 -3286 5226 -3234
rect 5174 -3376 5226 -3324
rect 5174 -3466 5226 -3414
rect 5174 -3556 5226 -3504
rect 5554 -3106 5606 -3054
rect 5554 -3196 5606 -3144
rect 5554 -3286 5606 -3234
rect 5554 -3376 5606 -3324
rect 5554 -3466 5606 -3414
rect 5554 -3556 5606 -3504
rect 5934 -3106 5986 -3054
rect 5934 -3196 5986 -3144
rect 5934 -3286 5986 -3234
rect 5934 -3376 5986 -3324
rect 5934 -3466 5986 -3414
rect 5934 -3556 5986 -3504
rect 6314 -3106 6366 -3054
rect 6314 -3196 6366 -3144
rect 6314 -3286 6366 -3234
rect 6314 -3376 6366 -3324
rect 6314 -3466 6366 -3414
rect 6314 -3556 6366 -3504
rect 6517 -2286 6569 -2234
rect 6581 -2286 6633 -2234
rect 6897 -2286 6949 -2234
rect 6961 -2286 7013 -2234
rect 7277 -2286 7329 -2234
rect 7341 -2286 7393 -2234
rect 7657 -2286 7709 -2234
rect 7721 -2286 7773 -2234
rect 8037 -2286 8089 -2234
rect 8101 -2286 8153 -2234
rect 6694 -3106 6746 -3054
rect 6694 -3196 6746 -3144
rect 6694 -3286 6746 -3234
rect 6694 -3376 6746 -3324
rect 6694 -3466 6746 -3414
rect 6694 -3556 6746 -3504
rect 7074 -3106 7126 -3054
rect 7074 -3196 7126 -3144
rect 7074 -3286 7126 -3234
rect 7074 -3376 7126 -3324
rect 7074 -3466 7126 -3414
rect 7074 -3556 7126 -3504
rect 7454 -3106 7506 -3054
rect 7454 -3196 7506 -3144
rect 7454 -3286 7506 -3234
rect 7454 -3376 7506 -3324
rect 7454 -3466 7506 -3414
rect 7454 -3556 7506 -3504
rect 7834 -3106 7886 -3054
rect 7834 -3196 7886 -3144
rect 7834 -3286 7886 -3234
rect 7834 -3376 7886 -3324
rect 7834 -3466 7886 -3414
rect 7834 -3556 7886 -3504
rect 8214 -3106 8266 -3054
rect 8214 -3196 8266 -3144
rect 8214 -3286 8266 -3234
rect 8214 -3376 8266 -3324
rect 8214 -3466 8266 -3414
rect 8214 -3556 8266 -3504
rect -236 -4346 -184 -4294
rect -236 -4736 -184 -4684
rect -236 -4816 -184 -4764
rect 437 -4346 489 -4294
rect 501 -4346 553 -4294
rect 817 -4346 869 -4294
rect 881 -4346 933 -4294
rect 1197 -4346 1249 -4294
rect 1261 -4346 1313 -4294
rect 1577 -4346 1629 -4294
rect 1641 -4346 1693 -4294
rect 1957 -4346 2009 -4294
rect 2021 -4346 2073 -4294
rect 2337 -4346 2389 -4294
rect 2401 -4346 2453 -4294
rect 2717 -4346 2769 -4294
rect 2781 -4346 2833 -4294
rect 3097 -4346 3149 -4294
rect 3161 -4346 3213 -4294
rect 3477 -4346 3529 -4294
rect 3541 -4346 3593 -4294
rect 3857 -4346 3909 -4294
rect 3921 -4346 3973 -4294
rect 4024 -4346 4076 -4294
rect 4124 -4346 4176 -4294
rect 4617 -4346 4669 -4294
rect 4681 -4346 4733 -4294
rect 4997 -4346 5049 -4294
rect 5061 -4346 5113 -4294
rect 5377 -4346 5429 -4294
rect 5441 -4346 5493 -4294
rect 5757 -4346 5809 -4294
rect 5821 -4346 5873 -4294
rect 6137 -4346 6189 -4294
rect 6201 -4346 6253 -4294
rect 6314 -4346 6366 -4294
rect 6404 -4346 6456 -4294
rect 6517 -4346 6569 -4294
rect 6581 -4346 6633 -4294
rect 6897 -4346 6949 -4294
rect 6961 -4346 7013 -4294
rect 7277 -4346 7329 -4294
rect 7341 -4346 7393 -4294
rect 7657 -4346 7709 -4294
rect 7721 -4346 7773 -4294
rect 8037 -4346 8089 -4294
rect 8101 -4346 8153 -4294
rect 8704 -2086 8756 -2034
rect 8704 -2166 8756 -2114
rect 8704 -4346 8756 -4294
rect 8704 -4426 8756 -4374
rect 8704 -5056 8756 -5004
rect 8704 -5136 8756 -5084
<< metal2 >>
rect 4470 5338 4570 5360
rect 4470 5282 4492 5338
rect 4548 5282 4570 5338
rect 4470 5100 4570 5282
rect -250 5088 8910 5100
rect -250 5032 -238 5088
rect -182 5032 -148 5088
rect -92 5086 8910 5088
rect -92 5034 8764 5086
rect 8816 5034 8844 5086
rect 8896 5034 8910 5086
rect -92 5032 8910 5034
rect -250 5020 8910 5032
rect 4160 4978 4570 4990
rect 4160 4922 4172 4978
rect 4228 4922 4262 4978
rect 4318 4922 4412 4978
rect 4468 4922 4502 4978
rect 4558 4922 4570 4978
rect 4160 4910 4570 4922
rect -110 4868 8770 4880
rect -110 4812 -98 4868
rect -42 4812 -8 4868
rect 48 4812 8612 4868
rect 8668 4812 8702 4868
rect 8758 4812 8770 4868
rect -110 4800 8770 4812
rect 220 4766 2290 4770
rect 220 4758 2144 4766
rect 220 4702 232 4758
rect 288 4702 322 4758
rect 378 4714 2144 4758
rect 2196 4714 2224 4766
rect 2276 4714 2290 4766
rect 378 4710 2290 4714
rect 378 4702 390 4710
rect 220 4690 390 4702
rect 1910 4426 2580 4430
rect 1910 4374 1934 4426
rect 1986 4374 2014 4426
rect 2066 4374 2334 4426
rect 2386 4374 2434 4426
rect 2486 4374 2580 4426
rect 1910 4370 2580 4374
rect -590 4310 -490 4350
rect 4130 4318 4330 4330
rect -590 4306 3990 4310
rect -590 4298 437 4306
rect -590 4250 -98 4298
rect -110 4242 -98 4250
rect -42 4254 437 4298
rect 489 4254 501 4306
rect 553 4254 817 4306
rect 869 4254 881 4306
rect 933 4254 1197 4306
rect 1249 4254 1261 4306
rect 1313 4254 1577 4306
rect 1629 4254 1641 4306
rect 1693 4254 1957 4306
rect 2009 4254 2021 4306
rect 2073 4254 2337 4306
rect 2389 4254 2401 4306
rect 2453 4254 2717 4306
rect 2769 4254 2781 4306
rect 2833 4254 3097 4306
rect 3149 4254 3161 4306
rect 3213 4254 3477 4306
rect 3529 4254 3541 4306
rect 3593 4254 3857 4306
rect 3909 4254 3921 4306
rect 3973 4254 3990 4306
rect -42 4250 3990 4254
rect 4130 4262 4172 4318
rect 4228 4262 4262 4318
rect 4318 4262 4330 4318
rect 4130 4250 4330 4262
rect 4490 4318 4700 4330
rect 4490 4262 4522 4318
rect 4578 4262 4612 4318
rect 4668 4310 4700 4318
rect 4668 4306 6270 4310
rect 4668 4262 4685 4306
rect 4490 4259 4614 4262
rect 4666 4259 4685 4262
rect 4490 4254 4685 4259
rect 4737 4254 4997 4306
rect 5049 4254 5061 4306
rect 5113 4254 5377 4306
rect 5429 4254 5441 4306
rect 5493 4254 5757 4306
rect 5809 4254 5821 4306
rect 5873 4254 6137 4306
rect 6189 4254 6201 4306
rect 6253 4254 6270 4306
rect 4490 4250 6270 4254
rect 6300 4250 6380 4310
rect 6500 4306 8910 4310
rect 6500 4254 6517 4306
rect 6569 4254 6581 4306
rect 6633 4254 6897 4306
rect 6949 4254 6961 4306
rect 7013 4254 7277 4306
rect 7329 4254 7341 4306
rect 7393 4254 7657 4306
rect 7709 4254 7721 4306
rect 7773 4254 8037 4306
rect 8089 4254 8101 4306
rect 8153 4254 8844 4306
rect 8896 4254 8910 4306
rect 6500 4250 8910 4254
rect -42 4242 -30 4250
rect -110 4208 -30 4242
rect -110 4152 -98 4208
rect -42 4152 -30 4208
rect -110 4140 -30 4152
rect 600 3528 680 3540
rect 600 3472 612 3528
rect 668 3472 680 3528
rect 600 3438 680 3472
rect 600 3382 612 3438
rect 668 3382 680 3438
rect 600 3348 680 3382
rect 600 3292 612 3348
rect 668 3292 680 3348
rect 600 3258 680 3292
rect 600 3202 612 3258
rect 668 3202 680 3258
rect 600 3168 680 3202
rect 600 3112 612 3168
rect 668 3112 680 3168
rect 600 3078 680 3112
rect 600 3022 612 3078
rect 668 3022 680 3078
rect 600 3010 680 3022
rect 980 3528 1060 3540
rect 980 3472 992 3528
rect 1048 3472 1060 3528
rect 980 3438 1060 3472
rect 980 3382 992 3438
rect 1048 3382 1060 3438
rect 980 3348 1060 3382
rect 980 3292 992 3348
rect 1048 3292 1060 3348
rect 980 3258 1060 3292
rect 980 3202 992 3258
rect 1048 3202 1060 3258
rect 980 3168 1060 3202
rect 980 3112 992 3168
rect 1048 3112 1060 3168
rect 980 3078 1060 3112
rect 980 3022 992 3078
rect 1048 3022 1060 3078
rect 980 3010 1060 3022
rect 1360 3528 1440 3540
rect 1360 3472 1372 3528
rect 1428 3472 1440 3528
rect 1360 3438 1440 3472
rect 1360 3382 1372 3438
rect 1428 3382 1440 3438
rect 1360 3348 1440 3382
rect 1360 3292 1372 3348
rect 1428 3292 1440 3348
rect 1360 3258 1440 3292
rect 1360 3202 1372 3258
rect 1428 3202 1440 3258
rect 1360 3168 1440 3202
rect 1360 3112 1372 3168
rect 1428 3112 1440 3168
rect 1360 3078 1440 3112
rect 1360 3022 1372 3078
rect 1428 3022 1440 3078
rect 1360 3010 1440 3022
rect 1740 3528 1820 3540
rect 1740 3472 1752 3528
rect 1808 3472 1820 3528
rect 1740 3438 1820 3472
rect 1740 3382 1752 3438
rect 1808 3382 1820 3438
rect 1740 3348 1820 3382
rect 1740 3292 1752 3348
rect 1808 3292 1820 3348
rect 1740 3258 1820 3292
rect 1740 3202 1752 3258
rect 1808 3202 1820 3258
rect 1740 3168 1820 3202
rect 1740 3112 1752 3168
rect 1808 3112 1820 3168
rect 1740 3078 1820 3112
rect 1740 3022 1752 3078
rect 1808 3022 1820 3078
rect 1740 3010 1820 3022
rect 2120 3528 2200 3540
rect 2120 3472 2132 3528
rect 2188 3472 2200 3528
rect 2120 3438 2200 3472
rect 2120 3382 2132 3438
rect 2188 3382 2200 3438
rect 2120 3348 2200 3382
rect 2120 3292 2132 3348
rect 2188 3292 2200 3348
rect 2120 3258 2200 3292
rect 2120 3202 2132 3258
rect 2188 3202 2200 3258
rect 2120 3168 2200 3202
rect 2120 3112 2132 3168
rect 2188 3112 2200 3168
rect 2120 3078 2200 3112
rect 2120 3022 2132 3078
rect 2188 3022 2200 3078
rect 2120 3010 2200 3022
rect 2500 3528 2580 3540
rect 2500 3472 2512 3528
rect 2568 3472 2580 3528
rect 2500 3438 2580 3472
rect 2500 3382 2512 3438
rect 2568 3382 2580 3438
rect 2500 3348 2580 3382
rect 2500 3292 2512 3348
rect 2568 3292 2580 3348
rect 2500 3258 2580 3292
rect 2500 3202 2512 3258
rect 2568 3202 2580 3258
rect 2500 3168 2580 3202
rect 2500 3112 2512 3168
rect 2568 3112 2580 3168
rect 2500 3078 2580 3112
rect 2500 3022 2512 3078
rect 2568 3022 2580 3078
rect 2500 3010 2580 3022
rect 2880 3528 2960 3540
rect 2880 3472 2892 3528
rect 2948 3472 2960 3528
rect 2880 3438 2960 3472
rect 2880 3382 2892 3438
rect 2948 3382 2960 3438
rect 2880 3348 2960 3382
rect 2880 3292 2892 3348
rect 2948 3292 2960 3348
rect 2880 3258 2960 3292
rect 2880 3202 2892 3258
rect 2948 3202 2960 3258
rect 2880 3168 2960 3202
rect 2880 3112 2892 3168
rect 2948 3112 2960 3168
rect 2880 3078 2960 3112
rect 2880 3022 2892 3078
rect 2948 3022 2960 3078
rect 2880 3010 2960 3022
rect 3260 3528 3340 3540
rect 3260 3472 3272 3528
rect 3328 3472 3340 3528
rect 3260 3438 3340 3472
rect 3260 3382 3272 3438
rect 3328 3382 3340 3438
rect 3260 3348 3340 3382
rect 3260 3292 3272 3348
rect 3328 3292 3340 3348
rect 3260 3258 3340 3292
rect 3260 3202 3272 3258
rect 3328 3202 3340 3258
rect 3260 3168 3340 3202
rect 3260 3112 3272 3168
rect 3328 3112 3340 3168
rect 3260 3078 3340 3112
rect 3260 3022 3272 3078
rect 3328 3022 3340 3078
rect 3260 3010 3340 3022
rect 3640 3528 3720 3540
rect 3640 3472 3652 3528
rect 3708 3472 3720 3528
rect 3640 3438 3720 3472
rect 3640 3382 3652 3438
rect 3708 3382 3720 3438
rect 3640 3348 3720 3382
rect 3640 3292 3652 3348
rect 3708 3292 3720 3348
rect 3640 3258 3720 3292
rect 3640 3202 3652 3258
rect 3708 3202 3720 3258
rect 3640 3168 3720 3202
rect 3640 3112 3652 3168
rect 3708 3112 3720 3168
rect 3640 3078 3720 3112
rect 3640 3022 3652 3078
rect 3708 3022 3720 3078
rect 3640 3010 3720 3022
rect 4020 3528 4100 3540
rect 4020 3472 4032 3528
rect 4088 3472 4100 3528
rect 4020 3438 4100 3472
rect 4020 3382 4032 3438
rect 4088 3382 4100 3438
rect 4020 3348 4100 3382
rect 4020 3292 4032 3348
rect 4088 3292 4100 3348
rect 4020 3258 4100 3292
rect 4020 3202 4032 3258
rect 4088 3202 4100 3258
rect 4020 3168 4100 3202
rect 4020 3112 4032 3168
rect 4088 3112 4100 3168
rect 4020 3078 4100 3112
rect 4020 3022 4032 3078
rect 4088 3022 4100 3078
rect 4020 3010 4100 3022
rect -110 2326 -30 2330
rect -110 2274 -96 2326
rect -44 2274 -30 2326
rect -110 2250 -30 2274
rect -110 2246 2090 2250
rect -110 2194 -96 2246
rect -44 2194 437 2246
rect 489 2194 501 2246
rect 553 2194 817 2246
rect 869 2194 881 2246
rect 933 2194 1197 2246
rect 1249 2194 1261 2246
rect 1313 2194 1577 2246
rect 1629 2194 1641 2246
rect 1693 2194 1957 2246
rect 2009 2194 2021 2246
rect 2073 2194 2090 2246
rect -110 2190 2090 2194
rect 2320 2246 3990 2250
rect 2320 2194 2337 2246
rect 2389 2194 2401 2246
rect 2453 2194 2717 2246
rect 2769 2194 2781 2246
rect 2833 2194 3097 2246
rect 3149 2194 3161 2246
rect 3213 2194 3477 2246
rect 3529 2194 3541 2246
rect 3593 2194 3857 2246
rect 3909 2194 3921 2246
rect 3973 2194 3990 2246
rect 2320 2190 3990 2194
rect -110 2126 3990 2130
rect -110 2118 437 2126
rect -110 2062 -98 2118
rect -42 2074 437 2118
rect 489 2074 501 2126
rect 553 2074 817 2126
rect 869 2074 881 2126
rect 933 2074 1197 2126
rect 1249 2074 1261 2126
rect 1313 2074 1577 2126
rect 1629 2074 1641 2126
rect 1693 2074 1957 2126
rect 2009 2074 2021 2126
rect 2073 2074 2337 2126
rect 2389 2074 2401 2126
rect 2453 2074 2717 2126
rect 2769 2074 2781 2126
rect 2833 2074 3097 2126
rect 3149 2074 3161 2126
rect 3213 2074 3477 2126
rect 3529 2074 3541 2126
rect 3593 2074 3857 2126
rect 3909 2074 3921 2126
rect 3973 2074 3990 2126
rect -42 2070 3990 2074
rect -42 2062 -30 2070
rect -110 2028 -30 2062
rect -110 1972 -98 2028
rect -42 1972 -30 2028
rect -110 1960 -30 1972
rect -110 1798 -30 1820
rect -110 1742 -98 1798
rect -42 1742 -30 1798
rect -110 1708 -30 1742
rect -110 1652 -98 1708
rect -42 1652 -30 1708
rect -110 1640 -30 1652
rect 600 1378 680 1390
rect 600 1322 612 1378
rect 668 1322 680 1378
rect 600 1288 680 1322
rect 600 1232 612 1288
rect 668 1232 680 1288
rect 600 1198 680 1232
rect 600 1142 612 1198
rect 668 1142 680 1198
rect 600 1108 680 1142
rect 600 1052 612 1108
rect 668 1052 680 1108
rect 600 1018 680 1052
rect 600 962 612 1018
rect 668 962 680 1018
rect 600 928 680 962
rect 600 872 612 928
rect 668 872 680 928
rect 600 860 680 872
rect 980 1378 1060 1390
rect 980 1322 992 1378
rect 1048 1322 1060 1378
rect 980 1288 1060 1322
rect 980 1232 992 1288
rect 1048 1232 1060 1288
rect 980 1198 1060 1232
rect 980 1142 992 1198
rect 1048 1142 1060 1198
rect 980 1108 1060 1142
rect 980 1052 992 1108
rect 1048 1052 1060 1108
rect 980 1018 1060 1052
rect 980 962 992 1018
rect 1048 962 1060 1018
rect 980 928 1060 962
rect 980 872 992 928
rect 1048 872 1060 928
rect 980 860 1060 872
rect 1360 1378 1440 1390
rect 1360 1322 1372 1378
rect 1428 1322 1440 1378
rect 1360 1288 1440 1322
rect 1360 1232 1372 1288
rect 1428 1232 1440 1288
rect 1360 1198 1440 1232
rect 1360 1142 1372 1198
rect 1428 1142 1440 1198
rect 1360 1108 1440 1142
rect 1360 1052 1372 1108
rect 1428 1052 1440 1108
rect 1360 1018 1440 1052
rect 1360 962 1372 1018
rect 1428 962 1440 1018
rect 1360 928 1440 962
rect 1360 872 1372 928
rect 1428 872 1440 928
rect 1360 860 1440 872
rect 1740 1378 1820 1390
rect 1740 1322 1752 1378
rect 1808 1322 1820 1378
rect 1740 1288 1820 1322
rect 1740 1232 1752 1288
rect 1808 1232 1820 1288
rect 1740 1198 1820 1232
rect 1740 1142 1752 1198
rect 1808 1142 1820 1198
rect 1740 1108 1820 1142
rect 1740 1052 1752 1108
rect 1808 1052 1820 1108
rect 1740 1018 1820 1052
rect 1740 962 1752 1018
rect 1808 962 1820 1018
rect 1740 928 1820 962
rect 1740 872 1752 928
rect 1808 872 1820 928
rect 1740 860 1820 872
rect 2120 1378 2200 1390
rect 2120 1322 2132 1378
rect 2188 1322 2200 1378
rect 2120 1288 2200 1322
rect 2120 1232 2132 1288
rect 2188 1232 2200 1288
rect 2120 1198 2200 1232
rect 2120 1142 2132 1198
rect 2188 1142 2200 1198
rect 2120 1108 2200 1142
rect 2120 1052 2132 1108
rect 2188 1052 2200 1108
rect 2120 1018 2200 1052
rect 2120 962 2132 1018
rect 2188 962 2200 1018
rect 2120 928 2200 962
rect 2120 872 2132 928
rect 2188 872 2200 928
rect 2120 860 2200 872
rect 2500 1378 2580 1390
rect 2500 1322 2512 1378
rect 2568 1322 2580 1378
rect 2500 1288 2580 1322
rect 2500 1232 2512 1288
rect 2568 1232 2580 1288
rect 2500 1198 2580 1232
rect 2500 1142 2512 1198
rect 2568 1142 2580 1198
rect 2500 1108 2580 1142
rect 2500 1052 2512 1108
rect 2568 1052 2580 1108
rect 2500 1018 2580 1052
rect 2500 962 2512 1018
rect 2568 962 2580 1018
rect 2500 928 2580 962
rect 2500 872 2512 928
rect 2568 872 2580 928
rect 2500 860 2580 872
rect 2880 1378 2960 1390
rect 2880 1322 2892 1378
rect 2948 1322 2960 1378
rect 2880 1288 2960 1322
rect 2880 1232 2892 1288
rect 2948 1232 2960 1288
rect 2880 1198 2960 1232
rect 2880 1142 2892 1198
rect 2948 1142 2960 1198
rect 2880 1108 2960 1142
rect 2880 1052 2892 1108
rect 2948 1052 2960 1108
rect 2880 1018 2960 1052
rect 2880 962 2892 1018
rect 2948 962 2960 1018
rect 2880 928 2960 962
rect 2880 872 2892 928
rect 2948 872 2960 928
rect 2880 860 2960 872
rect 3260 1378 3340 1390
rect 3260 1322 3272 1378
rect 3328 1322 3340 1378
rect 3260 1288 3340 1322
rect 3260 1232 3272 1288
rect 3328 1232 3340 1288
rect 3260 1198 3340 1232
rect 3260 1142 3272 1198
rect 3328 1142 3340 1198
rect 3260 1108 3340 1142
rect 3260 1052 3272 1108
rect 3328 1052 3340 1108
rect 3260 1018 3340 1052
rect 3260 962 3272 1018
rect 3328 962 3340 1018
rect 3260 928 3340 962
rect 3260 872 3272 928
rect 3328 872 3340 928
rect 3260 860 3340 872
rect 3640 1378 3720 1390
rect 3640 1322 3652 1378
rect 3708 1322 3720 1378
rect 3640 1288 3720 1322
rect 3640 1232 3652 1288
rect 3708 1232 3720 1288
rect 3640 1198 3720 1232
rect 3640 1142 3652 1198
rect 3708 1142 3720 1198
rect 3640 1108 3720 1142
rect 3640 1052 3652 1108
rect 3708 1052 3720 1108
rect 3640 1018 3720 1052
rect 3640 962 3652 1018
rect 3708 962 3720 1018
rect 3640 928 3720 962
rect 3640 872 3652 928
rect 3708 872 3720 928
rect 3640 860 3720 872
rect 4020 1378 4100 1390
rect 4020 1322 4032 1378
rect 4088 1322 4100 1378
rect 4020 1288 4100 1322
rect 4020 1232 4032 1288
rect 4088 1232 4100 1288
rect 4020 1198 4100 1232
rect 4020 1142 4032 1198
rect 4088 1142 4100 1198
rect 4020 1108 4100 1142
rect 4020 1052 4032 1108
rect 4088 1052 4100 1108
rect 4020 1018 4100 1052
rect 4020 962 4032 1018
rect 4088 962 4100 1018
rect 4020 928 4100 962
rect 4020 872 4032 928
rect 4088 872 4100 928
rect 4020 860 4100 872
rect -110 168 -30 180
rect -110 112 -98 168
rect -42 112 -30 168
rect -110 78 -30 112
rect -250 48 -170 60
rect -250 -8 -238 48
rect -182 -8 -170 48
rect -110 22 -98 78
rect -42 70 -30 78
rect -42 66 2090 70
rect -42 22 437 66
rect -110 14 437 22
rect 489 14 501 66
rect 553 14 817 66
rect 869 14 881 66
rect 933 14 1197 66
rect 1249 14 1261 66
rect 1313 14 1577 66
rect 1629 14 1641 66
rect 1693 14 1957 66
rect 2009 14 2021 66
rect 2073 14 2090 66
rect -110 10 2090 14
rect 2320 66 3990 70
rect 2320 14 2337 66
rect 2389 14 2401 66
rect 2453 14 2717 66
rect 2769 14 2781 66
rect 2833 14 3097 66
rect 3149 14 3161 66
rect 3213 14 3477 66
rect 3529 14 3541 66
rect 3593 14 3857 66
rect 3909 14 3921 66
rect 3973 14 3990 66
rect 2320 10 3990 14
rect -250 -42 -170 -8
rect -250 -98 -238 -42
rect -182 -50 -170 -42
rect 4130 -50 4190 4250
rect 8830 4226 8910 4250
rect 8830 4174 8844 4226
rect 8896 4174 8910 4226
rect 8830 4170 8910 4174
rect 4780 3528 4860 3540
rect 4780 3472 4792 3528
rect 4848 3472 4860 3528
rect 4780 3438 4860 3472
rect 4780 3382 4792 3438
rect 4848 3382 4860 3438
rect 4780 3348 4860 3382
rect 4780 3292 4792 3348
rect 4848 3292 4860 3348
rect 4780 3258 4860 3292
rect 4780 3202 4792 3258
rect 4848 3202 4860 3258
rect 4780 3168 4860 3202
rect 4780 3112 4792 3168
rect 4848 3112 4860 3168
rect 4780 3078 4860 3112
rect 4780 3022 4792 3078
rect 4848 3022 4860 3078
rect 4780 3010 4860 3022
rect 5160 3528 5240 3540
rect 5160 3472 5172 3528
rect 5228 3472 5240 3528
rect 5160 3438 5240 3472
rect 5160 3382 5172 3438
rect 5228 3382 5240 3438
rect 5160 3348 5240 3382
rect 5160 3292 5172 3348
rect 5228 3292 5240 3348
rect 5160 3258 5240 3292
rect 5160 3202 5172 3258
rect 5228 3202 5240 3258
rect 5160 3168 5240 3202
rect 5160 3112 5172 3168
rect 5228 3112 5240 3168
rect 5160 3078 5240 3112
rect 5160 3022 5172 3078
rect 5228 3022 5240 3078
rect 5160 3010 5240 3022
rect 5540 3528 5620 3540
rect 5540 3472 5552 3528
rect 5608 3472 5620 3528
rect 5540 3438 5620 3472
rect 5540 3382 5552 3438
rect 5608 3382 5620 3438
rect 5540 3348 5620 3382
rect 5540 3292 5552 3348
rect 5608 3292 5620 3348
rect 5540 3258 5620 3292
rect 5540 3202 5552 3258
rect 5608 3202 5620 3258
rect 5540 3168 5620 3202
rect 5540 3112 5552 3168
rect 5608 3112 5620 3168
rect 5540 3078 5620 3112
rect 5540 3022 5552 3078
rect 5608 3022 5620 3078
rect 5540 3010 5620 3022
rect 5920 3528 6000 3540
rect 5920 3472 5932 3528
rect 5988 3472 6000 3528
rect 5920 3438 6000 3472
rect 5920 3382 5932 3438
rect 5988 3382 6000 3438
rect 5920 3348 6000 3382
rect 5920 3292 5932 3348
rect 5988 3292 6000 3348
rect 5920 3258 6000 3292
rect 5920 3202 5932 3258
rect 5988 3202 6000 3258
rect 5920 3168 6000 3202
rect 5920 3112 5932 3168
rect 5988 3112 6000 3168
rect 5920 3078 6000 3112
rect 5920 3022 5932 3078
rect 5988 3022 6000 3078
rect 5920 3010 6000 3022
rect 6300 3528 6380 3540
rect 6300 3472 6312 3528
rect 6368 3472 6380 3528
rect 6300 3438 6380 3472
rect 6300 3382 6312 3438
rect 6368 3382 6380 3438
rect 6300 3348 6380 3382
rect 6300 3292 6312 3348
rect 6368 3292 6380 3348
rect 6300 3258 6380 3292
rect 6300 3202 6312 3258
rect 6368 3202 6380 3258
rect 6300 3168 6380 3202
rect 6300 3112 6312 3168
rect 6368 3112 6380 3168
rect 6300 3078 6380 3112
rect 6300 3022 6312 3078
rect 6368 3022 6380 3078
rect 6300 3010 6380 3022
rect 6680 3528 6760 3540
rect 6680 3472 6692 3528
rect 6748 3472 6760 3528
rect 6680 3438 6760 3472
rect 6680 3382 6692 3438
rect 6748 3382 6760 3438
rect 6680 3348 6760 3382
rect 6680 3292 6692 3348
rect 6748 3292 6760 3348
rect 6680 3258 6760 3292
rect 6680 3202 6692 3258
rect 6748 3202 6760 3258
rect 6680 3168 6760 3202
rect 6680 3112 6692 3168
rect 6748 3112 6760 3168
rect 6680 3078 6760 3112
rect 6680 3022 6692 3078
rect 6748 3022 6760 3078
rect 6680 3010 6760 3022
rect 7060 3528 7140 3540
rect 7060 3472 7072 3528
rect 7128 3472 7140 3528
rect 7060 3438 7140 3472
rect 7060 3382 7072 3438
rect 7128 3382 7140 3438
rect 7060 3348 7140 3382
rect 7060 3292 7072 3348
rect 7128 3292 7140 3348
rect 7060 3258 7140 3292
rect 7060 3202 7072 3258
rect 7128 3202 7140 3258
rect 7060 3168 7140 3202
rect 7060 3112 7072 3168
rect 7128 3112 7140 3168
rect 7060 3078 7140 3112
rect 7060 3022 7072 3078
rect 7128 3022 7140 3078
rect 7060 3010 7140 3022
rect 7440 3528 7520 3540
rect 7440 3472 7452 3528
rect 7508 3472 7520 3528
rect 7440 3438 7520 3472
rect 7440 3382 7452 3438
rect 7508 3382 7520 3438
rect 7440 3348 7520 3382
rect 7440 3292 7452 3348
rect 7508 3292 7520 3348
rect 7440 3258 7520 3292
rect 7440 3202 7452 3258
rect 7508 3202 7520 3258
rect 7440 3168 7520 3202
rect 7440 3112 7452 3168
rect 7508 3112 7520 3168
rect 7440 3078 7520 3112
rect 7440 3022 7452 3078
rect 7508 3022 7520 3078
rect 7440 3010 7520 3022
rect 7820 3528 7900 3540
rect 7820 3472 7832 3528
rect 7888 3472 7900 3528
rect 7820 3438 7900 3472
rect 7820 3382 7832 3438
rect 7888 3382 7900 3438
rect 7820 3348 7900 3382
rect 7820 3292 7832 3348
rect 7888 3292 7900 3348
rect 7820 3258 7900 3292
rect 7820 3202 7832 3258
rect 7888 3202 7900 3258
rect 7820 3168 7900 3202
rect 7820 3112 7832 3168
rect 7888 3112 7900 3168
rect 7820 3078 7900 3112
rect 7820 3022 7832 3078
rect 7888 3022 7900 3078
rect 7820 3010 7900 3022
rect 8200 3528 8280 3540
rect 8200 3472 8212 3528
rect 8268 3472 8280 3528
rect 8200 3438 8280 3472
rect 8200 3382 8212 3438
rect 8268 3382 8280 3438
rect 8200 3348 8280 3382
rect 8200 3292 8212 3348
rect 8268 3292 8280 3348
rect 8200 3258 8280 3292
rect 8200 3202 8212 3258
rect 8268 3202 8280 3258
rect 8200 3168 8280 3202
rect 8200 3112 8212 3168
rect 8268 3112 8280 3168
rect 8200 3078 8280 3112
rect 8200 3022 8212 3078
rect 8268 3022 8280 3078
rect 8200 3010 8280 3022
rect 4490 2348 4570 2360
rect 4490 2292 4502 2348
rect 4558 2292 4570 2348
rect 4490 2258 4570 2292
rect 4490 2202 4502 2258
rect 4558 2250 4570 2258
rect 8830 2348 8910 2370
rect 8830 2292 8842 2348
rect 8898 2292 8910 2348
rect 8830 2258 8910 2292
rect 8830 2250 8842 2258
rect 4558 2246 6270 2250
rect 4558 2202 4617 2246
rect 4490 2194 4617 2202
rect 4669 2194 4681 2246
rect 4733 2194 4997 2246
rect 5049 2194 5061 2246
rect 5113 2194 5377 2246
rect 5429 2194 5441 2246
rect 5493 2194 5757 2246
rect 5809 2194 5821 2246
rect 5873 2194 6137 2246
rect 6189 2194 6201 2246
rect 6253 2194 6270 2246
rect 4490 2190 6270 2194
rect 6500 2246 8842 2250
rect 6500 2194 6517 2246
rect 6569 2194 6581 2246
rect 6633 2194 6897 2246
rect 6949 2194 6961 2246
rect 7013 2194 7277 2246
rect 7329 2194 7341 2246
rect 7393 2194 7657 2246
rect 7709 2194 7721 2246
rect 7773 2194 8037 2246
rect 8089 2194 8101 2246
rect 8153 2202 8842 2246
rect 8898 2202 8910 2258
rect 8153 2194 8910 2202
rect 6500 2190 8910 2194
rect 4220 2138 4390 2150
rect 4220 2082 4232 2138
rect 4288 2082 4322 2138
rect 4378 2082 4390 2138
rect 4220 2070 4390 2082
rect 4600 2126 6270 2130
rect 4600 2074 4617 2126
rect 4669 2074 4681 2126
rect 4733 2074 4997 2126
rect 5049 2074 5061 2126
rect 5113 2074 5377 2126
rect 5429 2074 5441 2126
rect 5493 2074 5757 2126
rect 5809 2074 5821 2126
rect 5873 2074 6137 2126
rect 6189 2074 6201 2126
rect 6253 2074 6270 2126
rect 4600 2070 6270 2074
rect 6500 2126 8910 2130
rect 6500 2074 6517 2126
rect 6569 2074 6581 2126
rect 6633 2074 6897 2126
rect 6949 2074 6961 2126
rect 7013 2074 7277 2126
rect 7329 2074 7341 2126
rect 7393 2074 7657 2126
rect 7709 2074 7721 2126
rect 7773 2074 8037 2126
rect 8089 2074 8101 2126
rect 8153 2074 8844 2126
rect 8896 2074 8910 2126
rect 6500 2070 8910 2074
rect 8830 2046 8910 2070
rect 8830 1994 8844 2046
rect 8896 1994 8910 2046
rect 8830 1990 8910 1994
rect 4780 1378 4860 1390
rect 4780 1322 4792 1378
rect 4848 1322 4860 1378
rect 4780 1288 4860 1322
rect 4780 1232 4792 1288
rect 4848 1232 4860 1288
rect 4780 1198 4860 1232
rect 4780 1142 4792 1198
rect 4848 1142 4860 1198
rect 4780 1108 4860 1142
rect 4780 1052 4792 1108
rect 4848 1052 4860 1108
rect 4780 1018 4860 1052
rect 4780 962 4792 1018
rect 4848 962 4860 1018
rect 4780 928 4860 962
rect 4780 872 4792 928
rect 4848 872 4860 928
rect 4780 860 4860 872
rect 5160 1378 5240 1390
rect 5160 1322 5172 1378
rect 5228 1322 5240 1378
rect 5160 1288 5240 1322
rect 5160 1232 5172 1288
rect 5228 1232 5240 1288
rect 5160 1198 5240 1232
rect 5160 1142 5172 1198
rect 5228 1142 5240 1198
rect 5160 1108 5240 1142
rect 5160 1052 5172 1108
rect 5228 1052 5240 1108
rect 5160 1018 5240 1052
rect 5160 962 5172 1018
rect 5228 962 5240 1018
rect 5160 928 5240 962
rect 5160 872 5172 928
rect 5228 872 5240 928
rect 5160 860 5240 872
rect 5540 1378 5620 1390
rect 5540 1322 5552 1378
rect 5608 1322 5620 1378
rect 5540 1288 5620 1322
rect 5540 1232 5552 1288
rect 5608 1232 5620 1288
rect 5540 1198 5620 1232
rect 5540 1142 5552 1198
rect 5608 1142 5620 1198
rect 5540 1108 5620 1142
rect 5540 1052 5552 1108
rect 5608 1052 5620 1108
rect 5540 1018 5620 1052
rect 5540 962 5552 1018
rect 5608 962 5620 1018
rect 5540 928 5620 962
rect 5540 872 5552 928
rect 5608 872 5620 928
rect 5540 860 5620 872
rect 5920 1378 6000 1390
rect 5920 1322 5932 1378
rect 5988 1322 6000 1378
rect 5920 1288 6000 1322
rect 5920 1232 5932 1288
rect 5988 1232 6000 1288
rect 5920 1198 6000 1232
rect 5920 1142 5932 1198
rect 5988 1142 6000 1198
rect 5920 1108 6000 1142
rect 5920 1052 5932 1108
rect 5988 1052 6000 1108
rect 5920 1018 6000 1052
rect 5920 962 5932 1018
rect 5988 962 6000 1018
rect 5920 928 6000 962
rect 5920 872 5932 928
rect 5988 872 6000 928
rect 5920 860 6000 872
rect 6300 1378 6380 1390
rect 6300 1322 6312 1378
rect 6368 1322 6380 1378
rect 6300 1288 6380 1322
rect 6300 1232 6312 1288
rect 6368 1232 6380 1288
rect 6300 1198 6380 1232
rect 6300 1142 6312 1198
rect 6368 1142 6380 1198
rect 6300 1108 6380 1142
rect 6300 1052 6312 1108
rect 6368 1052 6380 1108
rect 6300 1018 6380 1052
rect 6300 962 6312 1018
rect 6368 962 6380 1018
rect 6300 928 6380 962
rect 6300 872 6312 928
rect 6368 872 6380 928
rect 6300 860 6380 872
rect 6680 1378 6760 1390
rect 6680 1322 6692 1378
rect 6748 1322 6760 1378
rect 6680 1288 6760 1322
rect 6680 1232 6692 1288
rect 6748 1232 6760 1288
rect 6680 1198 6760 1232
rect 6680 1142 6692 1198
rect 6748 1142 6760 1198
rect 6680 1108 6760 1142
rect 6680 1052 6692 1108
rect 6748 1052 6760 1108
rect 6680 1018 6760 1052
rect 6680 962 6692 1018
rect 6748 962 6760 1018
rect 6680 928 6760 962
rect 6680 872 6692 928
rect 6748 872 6760 928
rect 6680 860 6760 872
rect 7060 1378 7140 1390
rect 7060 1322 7072 1378
rect 7128 1322 7140 1378
rect 7060 1288 7140 1322
rect 7060 1232 7072 1288
rect 7128 1232 7140 1288
rect 7060 1198 7140 1232
rect 7060 1142 7072 1198
rect 7128 1142 7140 1198
rect 7060 1108 7140 1142
rect 7060 1052 7072 1108
rect 7128 1052 7140 1108
rect 7060 1018 7140 1052
rect 7060 962 7072 1018
rect 7128 962 7140 1018
rect 7060 928 7140 962
rect 7060 872 7072 928
rect 7128 872 7140 928
rect 7060 860 7140 872
rect 7440 1378 7520 1390
rect 7440 1322 7452 1378
rect 7508 1322 7520 1378
rect 7440 1288 7520 1322
rect 7440 1232 7452 1288
rect 7508 1232 7520 1288
rect 7440 1198 7520 1232
rect 7440 1142 7452 1198
rect 7508 1142 7520 1198
rect 7440 1108 7520 1142
rect 7440 1052 7452 1108
rect 7508 1052 7520 1108
rect 7440 1018 7520 1052
rect 7440 962 7452 1018
rect 7508 962 7520 1018
rect 7440 928 7520 962
rect 7440 872 7452 928
rect 7508 872 7520 928
rect 7440 860 7520 872
rect 7820 1378 7900 1390
rect 7820 1322 7832 1378
rect 7888 1322 7900 1378
rect 7820 1288 7900 1322
rect 7820 1232 7832 1288
rect 7888 1232 7900 1288
rect 7820 1198 7900 1232
rect 7820 1142 7832 1198
rect 7888 1142 7900 1198
rect 7820 1108 7900 1142
rect 7820 1052 7832 1108
rect 7888 1052 7900 1108
rect 7820 1018 7900 1052
rect 7820 962 7832 1018
rect 7888 962 7900 1018
rect 7820 928 7900 962
rect 7820 872 7832 928
rect 7888 872 7900 928
rect 7820 860 7900 872
rect 8200 1378 8280 1390
rect 8200 1322 8212 1378
rect 8268 1322 8280 1378
rect 8200 1288 8280 1322
rect 8200 1232 8212 1288
rect 8268 1232 8280 1288
rect 8200 1198 8280 1232
rect 8200 1142 8212 1198
rect 8268 1142 8280 1198
rect 8200 1108 8280 1142
rect 8200 1052 8212 1108
rect 8268 1052 8280 1108
rect 8200 1018 8280 1052
rect 8200 962 8212 1018
rect 8268 962 8280 1018
rect 8200 928 8280 962
rect 8200 872 8212 928
rect 8268 872 8280 928
rect 8200 860 8280 872
rect 4490 168 4570 180
rect 4490 112 4502 168
rect 4558 112 4570 168
rect 4490 78 4570 112
rect 4490 22 4502 78
rect 4558 70 4570 78
rect 8830 168 8910 180
rect 8830 112 8842 168
rect 8898 112 8910 168
rect 8830 78 8910 112
rect 8830 70 8842 78
rect 4558 66 6270 70
rect 4558 22 4617 66
rect 4490 14 4617 22
rect 4669 14 4681 66
rect 4733 14 4997 66
rect 5049 14 5061 66
rect 5113 14 5377 66
rect 5429 14 5441 66
rect 5493 14 5757 66
rect 5809 14 5821 66
rect 5873 14 6137 66
rect 6189 14 6201 66
rect 6253 14 6270 66
rect 4490 10 6270 14
rect 6500 66 8842 70
rect 6500 14 6517 66
rect 6569 14 6581 66
rect 6633 14 6897 66
rect 6949 14 6961 66
rect 7013 14 7277 66
rect 7329 14 7341 66
rect 7393 14 7657 66
rect 7709 14 7721 66
rect 7773 14 8037 66
rect 8089 14 8101 66
rect 8153 22 8842 66
rect 8898 22 8910 78
rect 8153 14 8910 22
rect 6500 10 8910 14
rect -182 -54 2090 -50
rect -182 -98 437 -54
rect -250 -106 437 -98
rect 489 -106 501 -54
rect 553 -106 817 -54
rect 869 -106 881 -54
rect 933 -106 1197 -54
rect 1249 -106 1261 -54
rect 1313 -106 1577 -54
rect 1629 -106 1641 -54
rect 1693 -106 1957 -54
rect 2009 -106 2021 -54
rect 2073 -106 2090 -54
rect -250 -110 2090 -106
rect 2320 -54 4190 -50
rect 2320 -106 2337 -54
rect 2389 -106 2401 -54
rect 2453 -106 2717 -54
rect 2769 -106 2781 -54
rect 2833 -106 3097 -54
rect 3149 -106 3161 -54
rect 3213 -106 3477 -54
rect 3529 -106 3541 -54
rect 3593 -106 3857 -54
rect 3909 -106 3921 -54
rect 3973 -106 4190 -54
rect 2320 -110 4190 -106
rect 4600 -54 8770 -50
rect 4600 -106 4617 -54
rect 4669 -106 4681 -54
rect 4733 -106 4997 -54
rect 5049 -106 5061 -54
rect 5113 -106 5377 -54
rect 5429 -106 5441 -54
rect 5493 -106 5757 -54
rect 5809 -106 5821 -54
rect 5873 -106 6137 -54
rect 6189 -106 6201 -54
rect 6253 -106 6517 -54
rect 6569 -106 6581 -54
rect 6633 -106 6897 -54
rect 6949 -106 6961 -54
rect 7013 -106 7277 -54
rect 7329 -106 7341 -54
rect 7393 -106 7657 -54
rect 7709 -106 7721 -54
rect 7773 -106 8037 -54
rect 8089 -106 8101 -54
rect 8153 -62 8770 -54
rect 8153 -106 8702 -62
rect 4600 -110 8702 -106
rect 600 -862 680 -850
rect 600 -918 612 -862
rect 668 -918 680 -862
rect 600 -952 680 -918
rect 600 -1008 612 -952
rect 668 -1008 680 -952
rect 600 -1042 680 -1008
rect 600 -1098 612 -1042
rect 668 -1098 680 -1042
rect 600 -1132 680 -1098
rect 600 -1188 612 -1132
rect 668 -1188 680 -1132
rect 600 -1222 680 -1188
rect 600 -1278 612 -1222
rect 668 -1278 680 -1222
rect 600 -1312 680 -1278
rect 600 -1368 612 -1312
rect 668 -1368 680 -1312
rect 600 -1380 680 -1368
rect 980 -862 1060 -850
rect 980 -918 992 -862
rect 1048 -918 1060 -862
rect 980 -952 1060 -918
rect 980 -1008 992 -952
rect 1048 -1008 1060 -952
rect 980 -1042 1060 -1008
rect 980 -1098 992 -1042
rect 1048 -1098 1060 -1042
rect 980 -1132 1060 -1098
rect 980 -1188 992 -1132
rect 1048 -1188 1060 -1132
rect 980 -1222 1060 -1188
rect 980 -1278 992 -1222
rect 1048 -1278 1060 -1222
rect 980 -1312 1060 -1278
rect 980 -1368 992 -1312
rect 1048 -1368 1060 -1312
rect 980 -1380 1060 -1368
rect 1360 -862 1440 -850
rect 1360 -918 1372 -862
rect 1428 -918 1440 -862
rect 1360 -952 1440 -918
rect 1360 -1008 1372 -952
rect 1428 -1008 1440 -952
rect 1360 -1042 1440 -1008
rect 1360 -1098 1372 -1042
rect 1428 -1098 1440 -1042
rect 1360 -1132 1440 -1098
rect 1360 -1188 1372 -1132
rect 1428 -1188 1440 -1132
rect 1360 -1222 1440 -1188
rect 1360 -1278 1372 -1222
rect 1428 -1278 1440 -1222
rect 1360 -1312 1440 -1278
rect 1360 -1368 1372 -1312
rect 1428 -1368 1440 -1312
rect 1360 -1380 1440 -1368
rect 1740 -862 1820 -850
rect 1740 -918 1752 -862
rect 1808 -918 1820 -862
rect 1740 -952 1820 -918
rect 1740 -1008 1752 -952
rect 1808 -1008 1820 -952
rect 1740 -1042 1820 -1008
rect 1740 -1098 1752 -1042
rect 1808 -1098 1820 -1042
rect 1740 -1132 1820 -1098
rect 1740 -1188 1752 -1132
rect 1808 -1188 1820 -1132
rect 1740 -1222 1820 -1188
rect 1740 -1278 1752 -1222
rect 1808 -1278 1820 -1222
rect 1740 -1312 1820 -1278
rect 1740 -1368 1752 -1312
rect 1808 -1368 1820 -1312
rect 1740 -1380 1820 -1368
rect 2120 -862 2200 -850
rect 2120 -918 2132 -862
rect 2188 -918 2200 -862
rect 2120 -952 2200 -918
rect 2120 -1008 2132 -952
rect 2188 -1008 2200 -952
rect 2120 -1042 2200 -1008
rect 2120 -1098 2132 -1042
rect 2188 -1098 2200 -1042
rect 2120 -1132 2200 -1098
rect 2120 -1188 2132 -1132
rect 2188 -1188 2200 -1132
rect 2120 -1222 2200 -1188
rect 2120 -1278 2132 -1222
rect 2188 -1278 2200 -1222
rect 2120 -1312 2200 -1278
rect 2120 -1368 2132 -1312
rect 2188 -1368 2200 -1312
rect 2120 -1380 2200 -1368
rect 2500 -862 2580 -850
rect 2500 -918 2512 -862
rect 2568 -918 2580 -862
rect 2500 -952 2580 -918
rect 2500 -1008 2512 -952
rect 2568 -1008 2580 -952
rect 2500 -1042 2580 -1008
rect 2500 -1098 2512 -1042
rect 2568 -1098 2580 -1042
rect 2500 -1132 2580 -1098
rect 2500 -1188 2512 -1132
rect 2568 -1188 2580 -1132
rect 2500 -1222 2580 -1188
rect 2500 -1278 2512 -1222
rect 2568 -1278 2580 -1222
rect 2500 -1312 2580 -1278
rect 2500 -1368 2512 -1312
rect 2568 -1368 2580 -1312
rect 2500 -1380 2580 -1368
rect 2880 -862 2960 -850
rect 2880 -918 2892 -862
rect 2948 -918 2960 -862
rect 2880 -952 2960 -918
rect 2880 -1008 2892 -952
rect 2948 -1008 2960 -952
rect 2880 -1042 2960 -1008
rect 2880 -1098 2892 -1042
rect 2948 -1098 2960 -1042
rect 2880 -1132 2960 -1098
rect 2880 -1188 2892 -1132
rect 2948 -1188 2960 -1132
rect 2880 -1222 2960 -1188
rect 2880 -1278 2892 -1222
rect 2948 -1278 2960 -1222
rect 2880 -1312 2960 -1278
rect 2880 -1368 2892 -1312
rect 2948 -1368 2960 -1312
rect 2880 -1380 2960 -1368
rect 3260 -862 3340 -850
rect 3260 -918 3272 -862
rect 3328 -918 3340 -862
rect 3260 -952 3340 -918
rect 3260 -1008 3272 -952
rect 3328 -1008 3340 -952
rect 3260 -1042 3340 -1008
rect 3260 -1098 3272 -1042
rect 3328 -1098 3340 -1042
rect 3260 -1132 3340 -1098
rect 3260 -1188 3272 -1132
rect 3328 -1188 3340 -1132
rect 3260 -1222 3340 -1188
rect 3260 -1278 3272 -1222
rect 3328 -1278 3340 -1222
rect 3260 -1312 3340 -1278
rect 3260 -1368 3272 -1312
rect 3328 -1368 3340 -1312
rect 3260 -1380 3340 -1368
rect 3640 -862 3720 -850
rect 3640 -918 3652 -862
rect 3708 -918 3720 -862
rect 3640 -952 3720 -918
rect 3640 -1008 3652 -952
rect 3708 -1008 3720 -952
rect 3640 -1042 3720 -1008
rect 3640 -1098 3652 -1042
rect 3708 -1098 3720 -1042
rect 3640 -1132 3720 -1098
rect 3640 -1188 3652 -1132
rect 3708 -1188 3720 -1132
rect 3640 -1222 3720 -1188
rect 3640 -1278 3652 -1222
rect 3708 -1278 3720 -1222
rect 3640 -1312 3720 -1278
rect 3640 -1368 3652 -1312
rect 3708 -1368 3720 -1312
rect 3640 -1380 3720 -1368
rect 4020 -862 4100 -850
rect 4020 -918 4032 -862
rect 4088 -918 4100 -862
rect 4020 -952 4100 -918
rect 4020 -1008 4032 -952
rect 4088 -1008 4100 -952
rect 4020 -1042 4100 -1008
rect 4020 -1098 4032 -1042
rect 4088 -1098 4100 -1042
rect 4020 -1132 4100 -1098
rect 4020 -1188 4032 -1132
rect 4088 -1188 4100 -1132
rect 4020 -1222 4100 -1188
rect 4020 -1278 4032 -1222
rect 4088 -1278 4100 -1222
rect 4020 -1312 4100 -1278
rect 4020 -1368 4032 -1312
rect 4088 -1368 4100 -1312
rect 4020 -1380 4100 -1368
rect -250 -2034 -170 -2030
rect -250 -2086 -236 -2034
rect -184 -2086 -170 -2034
rect -590 -2110 -490 -2090
rect -250 -2110 -170 -2086
rect -590 -2112 2090 -2110
rect -590 -2168 -568 -2112
rect -512 -2114 2090 -2112
rect -512 -2166 -236 -2114
rect -184 -2166 437 -2114
rect 489 -2166 501 -2114
rect 553 -2166 817 -2114
rect 869 -2166 881 -2114
rect 933 -2166 1197 -2114
rect 1249 -2166 1261 -2114
rect 1313 -2166 1577 -2114
rect 1629 -2166 1641 -2114
rect 1693 -2166 1957 -2114
rect 2009 -2166 2021 -2114
rect 2073 -2166 2090 -2114
rect -512 -2168 2090 -2166
rect -590 -2170 2090 -2168
rect 2320 -2114 4070 -2110
rect 2320 -2166 2337 -2114
rect 2389 -2166 2401 -2114
rect 2453 -2166 2717 -2114
rect 2769 -2166 2781 -2114
rect 2833 -2166 3097 -2114
rect 3149 -2166 3161 -2114
rect 3213 -2166 3477 -2114
rect 3529 -2166 3541 -2114
rect 3593 -2166 3857 -2114
rect 3909 -2166 3921 -2114
rect 3973 -2166 4004 -2114
rect 4056 -2166 4070 -2114
rect 2320 -2170 4070 -2166
rect -590 -2190 -490 -2170
rect 4130 -2230 4190 -110
rect 8690 -118 8702 -110
rect 8758 -118 8770 -62
rect 8690 -152 8770 -118
rect 8690 -208 8702 -152
rect 8758 -208 8770 -152
rect 8690 -220 8770 -208
rect 4780 -862 4860 -850
rect 4780 -918 4792 -862
rect 4848 -918 4860 -862
rect 4780 -952 4860 -918
rect 4780 -1008 4792 -952
rect 4848 -1008 4860 -952
rect 4780 -1042 4860 -1008
rect 4780 -1098 4792 -1042
rect 4848 -1098 4860 -1042
rect 4780 -1132 4860 -1098
rect 4780 -1188 4792 -1132
rect 4848 -1188 4860 -1132
rect 4780 -1222 4860 -1188
rect 4780 -1278 4792 -1222
rect 4848 -1278 4860 -1222
rect 4780 -1312 4860 -1278
rect 4780 -1368 4792 -1312
rect 4848 -1368 4860 -1312
rect 4780 -1380 4860 -1368
rect 5160 -862 5240 -850
rect 5160 -918 5172 -862
rect 5228 -918 5240 -862
rect 5160 -952 5240 -918
rect 5160 -1008 5172 -952
rect 5228 -1008 5240 -952
rect 5160 -1042 5240 -1008
rect 5160 -1098 5172 -1042
rect 5228 -1098 5240 -1042
rect 5160 -1132 5240 -1098
rect 5160 -1188 5172 -1132
rect 5228 -1188 5240 -1132
rect 5160 -1222 5240 -1188
rect 5160 -1278 5172 -1222
rect 5228 -1278 5240 -1222
rect 5160 -1312 5240 -1278
rect 5160 -1368 5172 -1312
rect 5228 -1368 5240 -1312
rect 5160 -1380 5240 -1368
rect 5540 -862 5620 -850
rect 5540 -918 5552 -862
rect 5608 -918 5620 -862
rect 5540 -952 5620 -918
rect 5540 -1008 5552 -952
rect 5608 -1008 5620 -952
rect 5540 -1042 5620 -1008
rect 5540 -1098 5552 -1042
rect 5608 -1098 5620 -1042
rect 5540 -1132 5620 -1098
rect 5540 -1188 5552 -1132
rect 5608 -1188 5620 -1132
rect 5540 -1222 5620 -1188
rect 5540 -1278 5552 -1222
rect 5608 -1278 5620 -1222
rect 5540 -1312 5620 -1278
rect 5540 -1368 5552 -1312
rect 5608 -1368 5620 -1312
rect 5540 -1380 5620 -1368
rect 5920 -862 6000 -850
rect 5920 -918 5932 -862
rect 5988 -918 6000 -862
rect 5920 -952 6000 -918
rect 5920 -1008 5932 -952
rect 5988 -1008 6000 -952
rect 5920 -1042 6000 -1008
rect 5920 -1098 5932 -1042
rect 5988 -1098 6000 -1042
rect 5920 -1132 6000 -1098
rect 5920 -1188 5932 -1132
rect 5988 -1188 6000 -1132
rect 5920 -1222 6000 -1188
rect 5920 -1278 5932 -1222
rect 5988 -1278 6000 -1222
rect 5920 -1312 6000 -1278
rect 5920 -1368 5932 -1312
rect 5988 -1368 6000 -1312
rect 5920 -1380 6000 -1368
rect 6300 -862 6380 -850
rect 6300 -918 6312 -862
rect 6368 -918 6380 -862
rect 6300 -952 6380 -918
rect 6300 -1008 6312 -952
rect 6368 -1008 6380 -952
rect 6300 -1042 6380 -1008
rect 6300 -1098 6312 -1042
rect 6368 -1098 6380 -1042
rect 6300 -1132 6380 -1098
rect 6300 -1188 6312 -1132
rect 6368 -1188 6380 -1132
rect 6300 -1222 6380 -1188
rect 6300 -1278 6312 -1222
rect 6368 -1278 6380 -1222
rect 6300 -1312 6380 -1278
rect 6300 -1368 6312 -1312
rect 6368 -1368 6380 -1312
rect 6300 -1380 6380 -1368
rect 6680 -862 6760 -850
rect 6680 -918 6692 -862
rect 6748 -918 6760 -862
rect 6680 -952 6760 -918
rect 6680 -1008 6692 -952
rect 6748 -1008 6760 -952
rect 6680 -1042 6760 -1008
rect 6680 -1098 6692 -1042
rect 6748 -1098 6760 -1042
rect 6680 -1132 6760 -1098
rect 6680 -1188 6692 -1132
rect 6748 -1188 6760 -1132
rect 6680 -1222 6760 -1188
rect 6680 -1278 6692 -1222
rect 6748 -1278 6760 -1222
rect 6680 -1312 6760 -1278
rect 6680 -1368 6692 -1312
rect 6748 -1368 6760 -1312
rect 6680 -1380 6760 -1368
rect 7060 -862 7140 -850
rect 7060 -918 7072 -862
rect 7128 -918 7140 -862
rect 7060 -952 7140 -918
rect 7060 -1008 7072 -952
rect 7128 -1008 7140 -952
rect 7060 -1042 7140 -1008
rect 7060 -1098 7072 -1042
rect 7128 -1098 7140 -1042
rect 7060 -1132 7140 -1098
rect 7060 -1188 7072 -1132
rect 7128 -1188 7140 -1132
rect 7060 -1222 7140 -1188
rect 7060 -1278 7072 -1222
rect 7128 -1278 7140 -1222
rect 7060 -1312 7140 -1278
rect 7060 -1368 7072 -1312
rect 7128 -1368 7140 -1312
rect 7060 -1380 7140 -1368
rect 7440 -862 7520 -850
rect 7440 -918 7452 -862
rect 7508 -918 7520 -862
rect 7440 -952 7520 -918
rect 7440 -1008 7452 -952
rect 7508 -1008 7520 -952
rect 7440 -1042 7520 -1008
rect 7440 -1098 7452 -1042
rect 7508 -1098 7520 -1042
rect 7440 -1132 7520 -1098
rect 7440 -1188 7452 -1132
rect 7508 -1188 7520 -1132
rect 7440 -1222 7520 -1188
rect 7440 -1278 7452 -1222
rect 7508 -1278 7520 -1222
rect 7440 -1312 7520 -1278
rect 7440 -1368 7452 -1312
rect 7508 -1368 7520 -1312
rect 7440 -1380 7520 -1368
rect 7820 -862 7900 -850
rect 7820 -918 7832 -862
rect 7888 -918 7900 -862
rect 7820 -952 7900 -918
rect 7820 -1008 7832 -952
rect 7888 -1008 7900 -952
rect 7820 -1042 7900 -1008
rect 7820 -1098 7832 -1042
rect 7888 -1098 7900 -1042
rect 7820 -1132 7900 -1098
rect 7820 -1188 7832 -1132
rect 7888 -1188 7900 -1132
rect 7820 -1222 7900 -1188
rect 7820 -1278 7832 -1222
rect 7888 -1278 7900 -1222
rect 7820 -1312 7900 -1278
rect 7820 -1368 7832 -1312
rect 7888 -1368 7900 -1312
rect 7820 -1380 7900 -1368
rect 8200 -862 8280 -850
rect 8200 -918 8212 -862
rect 8268 -918 8280 -862
rect 8200 -952 8280 -918
rect 8200 -1008 8212 -952
rect 8268 -1008 8280 -952
rect 8200 -1042 8280 -1008
rect 8200 -1098 8212 -1042
rect 8268 -1098 8280 -1042
rect 8200 -1132 8280 -1098
rect 8200 -1188 8212 -1132
rect 8268 -1188 8280 -1132
rect 8200 -1222 8280 -1188
rect 8200 -1278 8212 -1222
rect 8268 -1278 8280 -1222
rect 8200 -1312 8280 -1278
rect 8200 -1368 8212 -1312
rect 8268 -1368 8280 -1312
rect 8200 -1380 8280 -1368
rect 8690 -2034 8770 -2030
rect 8690 -2086 8704 -2034
rect 8756 -2086 8770 -2034
rect 8690 -2110 8770 -2086
rect 4600 -2114 6270 -2110
rect 4600 -2166 4617 -2114
rect 4669 -2166 4681 -2114
rect 4733 -2166 4997 -2114
rect 5049 -2166 5061 -2114
rect 5113 -2166 5377 -2114
rect 5429 -2166 5441 -2114
rect 5493 -2166 5757 -2114
rect 5809 -2166 5821 -2114
rect 5873 -2166 6137 -2114
rect 6189 -2166 6201 -2114
rect 6253 -2166 6270 -2114
rect 4600 -2170 6270 -2166
rect 6500 -2114 8770 -2110
rect 6500 -2166 6517 -2114
rect 6569 -2166 6581 -2114
rect 6633 -2166 6897 -2114
rect 6949 -2166 6961 -2114
rect 7013 -2166 7277 -2114
rect 7329 -2166 7341 -2114
rect 7393 -2166 7657 -2114
rect 7709 -2166 7721 -2114
rect 7773 -2166 8037 -2114
rect 8089 -2166 8101 -2114
rect 8153 -2166 8704 -2114
rect 8756 -2166 8770 -2114
rect 6500 -2170 8770 -2166
rect -250 -2234 2090 -2230
rect -250 -2242 437 -2234
rect -250 -2298 -238 -2242
rect -182 -2286 437 -2242
rect 489 -2286 501 -2234
rect 553 -2286 817 -2234
rect 869 -2286 881 -2234
rect 933 -2286 1197 -2234
rect 1249 -2286 1261 -2234
rect 1313 -2286 1577 -2234
rect 1629 -2286 1641 -2234
rect 1693 -2286 1957 -2234
rect 2009 -2286 2021 -2234
rect 2073 -2286 2090 -2234
rect -182 -2290 2090 -2286
rect 2320 -2234 4190 -2230
rect 2320 -2286 2337 -2234
rect 2389 -2286 2401 -2234
rect 2453 -2286 2717 -2234
rect 2769 -2286 2781 -2234
rect 2833 -2286 3097 -2234
rect 3149 -2286 3161 -2234
rect 3213 -2286 3477 -2234
rect 3529 -2286 3541 -2234
rect 3593 -2286 3857 -2234
rect 3909 -2286 3921 -2234
rect 3973 -2286 4190 -2234
rect 2320 -2290 4190 -2286
rect 4600 -2234 8770 -2230
rect 4600 -2286 4617 -2234
rect 4669 -2286 4681 -2234
rect 4733 -2286 4997 -2234
rect 5049 -2286 5061 -2234
rect 5113 -2286 5377 -2234
rect 5429 -2286 5441 -2234
rect 5493 -2286 5757 -2234
rect 5809 -2286 5821 -2234
rect 5873 -2286 6137 -2234
rect 6189 -2286 6201 -2234
rect 6253 -2286 6517 -2234
rect 6569 -2286 6581 -2234
rect 6633 -2286 6897 -2234
rect 6949 -2286 6961 -2234
rect 7013 -2286 7277 -2234
rect 7329 -2286 7341 -2234
rect 7393 -2286 7657 -2234
rect 7709 -2286 7721 -2234
rect 7773 -2286 8037 -2234
rect 8089 -2286 8101 -2234
rect 8153 -2242 8770 -2234
rect 8153 -2286 8702 -2242
rect 4600 -2290 8702 -2286
rect -182 -2298 -170 -2290
rect -250 -2332 -170 -2298
rect -250 -2388 -238 -2332
rect -182 -2388 -170 -2332
rect -250 -2400 -170 -2388
rect 8690 -2298 8702 -2290
rect 8758 -2298 8770 -2242
rect 8690 -2332 8770 -2298
rect 8690 -2388 8702 -2332
rect 8758 -2388 8770 -2332
rect 8690 -2400 8770 -2388
rect 600 -3052 680 -3040
rect 600 -3108 612 -3052
rect 668 -3108 680 -3052
rect 600 -3142 680 -3108
rect 600 -3198 612 -3142
rect 668 -3198 680 -3142
rect 600 -3232 680 -3198
rect 600 -3288 612 -3232
rect 668 -3288 680 -3232
rect 600 -3322 680 -3288
rect 600 -3378 612 -3322
rect 668 -3378 680 -3322
rect 600 -3412 680 -3378
rect 600 -3468 612 -3412
rect 668 -3468 680 -3412
rect 600 -3502 680 -3468
rect 600 -3558 612 -3502
rect 668 -3558 680 -3502
rect 600 -3570 680 -3558
rect 980 -3052 1060 -3040
rect 980 -3108 992 -3052
rect 1048 -3108 1060 -3052
rect 980 -3142 1060 -3108
rect 980 -3198 992 -3142
rect 1048 -3198 1060 -3142
rect 980 -3232 1060 -3198
rect 980 -3288 992 -3232
rect 1048 -3288 1060 -3232
rect 980 -3322 1060 -3288
rect 980 -3378 992 -3322
rect 1048 -3378 1060 -3322
rect 980 -3412 1060 -3378
rect 980 -3468 992 -3412
rect 1048 -3468 1060 -3412
rect 980 -3502 1060 -3468
rect 980 -3558 992 -3502
rect 1048 -3558 1060 -3502
rect 980 -3570 1060 -3558
rect 1360 -3052 1440 -3040
rect 1360 -3108 1372 -3052
rect 1428 -3108 1440 -3052
rect 1360 -3142 1440 -3108
rect 1360 -3198 1372 -3142
rect 1428 -3198 1440 -3142
rect 1360 -3232 1440 -3198
rect 1360 -3288 1372 -3232
rect 1428 -3288 1440 -3232
rect 1360 -3322 1440 -3288
rect 1360 -3378 1372 -3322
rect 1428 -3378 1440 -3322
rect 1360 -3412 1440 -3378
rect 1360 -3468 1372 -3412
rect 1428 -3468 1440 -3412
rect 1360 -3502 1440 -3468
rect 1360 -3558 1372 -3502
rect 1428 -3558 1440 -3502
rect 1360 -3570 1440 -3558
rect 1740 -3052 1820 -3040
rect 1740 -3108 1752 -3052
rect 1808 -3108 1820 -3052
rect 1740 -3142 1820 -3108
rect 1740 -3198 1752 -3142
rect 1808 -3198 1820 -3142
rect 1740 -3232 1820 -3198
rect 1740 -3288 1752 -3232
rect 1808 -3288 1820 -3232
rect 1740 -3322 1820 -3288
rect 1740 -3378 1752 -3322
rect 1808 -3378 1820 -3322
rect 1740 -3412 1820 -3378
rect 1740 -3468 1752 -3412
rect 1808 -3468 1820 -3412
rect 1740 -3502 1820 -3468
rect 1740 -3558 1752 -3502
rect 1808 -3558 1820 -3502
rect 1740 -3570 1820 -3558
rect 2120 -3052 2200 -3040
rect 2120 -3108 2132 -3052
rect 2188 -3108 2200 -3052
rect 2120 -3142 2200 -3108
rect 2120 -3198 2132 -3142
rect 2188 -3198 2200 -3142
rect 2120 -3232 2200 -3198
rect 2120 -3288 2132 -3232
rect 2188 -3288 2200 -3232
rect 2120 -3322 2200 -3288
rect 2120 -3378 2132 -3322
rect 2188 -3378 2200 -3322
rect 2120 -3412 2200 -3378
rect 2120 -3468 2132 -3412
rect 2188 -3468 2200 -3412
rect 2120 -3502 2200 -3468
rect 2120 -3558 2132 -3502
rect 2188 -3558 2200 -3502
rect 2120 -3570 2200 -3558
rect 2500 -3052 2580 -3040
rect 2500 -3108 2512 -3052
rect 2568 -3108 2580 -3052
rect 2500 -3142 2580 -3108
rect 2500 -3198 2512 -3142
rect 2568 -3198 2580 -3142
rect 2500 -3232 2580 -3198
rect 2500 -3288 2512 -3232
rect 2568 -3288 2580 -3232
rect 2500 -3322 2580 -3288
rect 2500 -3378 2512 -3322
rect 2568 -3378 2580 -3322
rect 2500 -3412 2580 -3378
rect 2500 -3468 2512 -3412
rect 2568 -3468 2580 -3412
rect 2500 -3502 2580 -3468
rect 2500 -3558 2512 -3502
rect 2568 -3558 2580 -3502
rect 2500 -3570 2580 -3558
rect 2880 -3052 2960 -3040
rect 2880 -3108 2892 -3052
rect 2948 -3108 2960 -3052
rect 2880 -3142 2960 -3108
rect 2880 -3198 2892 -3142
rect 2948 -3198 2960 -3142
rect 2880 -3232 2960 -3198
rect 2880 -3288 2892 -3232
rect 2948 -3288 2960 -3232
rect 2880 -3322 2960 -3288
rect 2880 -3378 2892 -3322
rect 2948 -3378 2960 -3322
rect 2880 -3412 2960 -3378
rect 2880 -3468 2892 -3412
rect 2948 -3468 2960 -3412
rect 2880 -3502 2960 -3468
rect 2880 -3558 2892 -3502
rect 2948 -3558 2960 -3502
rect 2880 -3570 2960 -3558
rect 3260 -3052 3340 -3040
rect 3260 -3108 3272 -3052
rect 3328 -3108 3340 -3052
rect 3260 -3142 3340 -3108
rect 3260 -3198 3272 -3142
rect 3328 -3198 3340 -3142
rect 3260 -3232 3340 -3198
rect 3260 -3288 3272 -3232
rect 3328 -3288 3340 -3232
rect 3260 -3322 3340 -3288
rect 3260 -3378 3272 -3322
rect 3328 -3378 3340 -3322
rect 3260 -3412 3340 -3378
rect 3260 -3468 3272 -3412
rect 3328 -3468 3340 -3412
rect 3260 -3502 3340 -3468
rect 3260 -3558 3272 -3502
rect 3328 -3558 3340 -3502
rect 3260 -3570 3340 -3558
rect 3640 -3052 3720 -3040
rect 3640 -3108 3652 -3052
rect 3708 -3108 3720 -3052
rect 3640 -3142 3720 -3108
rect 3640 -3198 3652 -3142
rect 3708 -3198 3720 -3142
rect 3640 -3232 3720 -3198
rect 3640 -3288 3652 -3232
rect 3708 -3288 3720 -3232
rect 3640 -3322 3720 -3288
rect 3640 -3378 3652 -3322
rect 3708 -3378 3720 -3322
rect 3640 -3412 3720 -3378
rect 3640 -3468 3652 -3412
rect 3708 -3468 3720 -3412
rect 3640 -3502 3720 -3468
rect 3640 -3558 3652 -3502
rect 3708 -3558 3720 -3502
rect 3640 -3570 3720 -3558
rect 4020 -3052 4100 -3040
rect 4020 -3108 4032 -3052
rect 4088 -3108 4100 -3052
rect 4020 -3142 4100 -3108
rect 4020 -3198 4032 -3142
rect 4088 -3198 4100 -3142
rect 4020 -3232 4100 -3198
rect 4020 -3288 4032 -3232
rect 4088 -3288 4100 -3232
rect 4020 -3322 4100 -3288
rect 4020 -3378 4032 -3322
rect 4088 -3378 4100 -3322
rect 4020 -3412 4100 -3378
rect 4020 -3468 4032 -3412
rect 4088 -3468 4100 -3412
rect 4020 -3502 4100 -3468
rect 4020 -3558 4032 -3502
rect 4088 -3558 4100 -3502
rect 4020 -3570 4100 -3558
rect 4780 -3052 4860 -3040
rect 4780 -3108 4792 -3052
rect 4848 -3108 4860 -3052
rect 4780 -3142 4860 -3108
rect 4780 -3198 4792 -3142
rect 4848 -3198 4860 -3142
rect 4780 -3232 4860 -3198
rect 4780 -3288 4792 -3232
rect 4848 -3288 4860 -3232
rect 4780 -3322 4860 -3288
rect 4780 -3378 4792 -3322
rect 4848 -3378 4860 -3322
rect 4780 -3412 4860 -3378
rect 4780 -3468 4792 -3412
rect 4848 -3468 4860 -3412
rect 4780 -3502 4860 -3468
rect 4780 -3558 4792 -3502
rect 4848 -3558 4860 -3502
rect 4780 -3570 4860 -3558
rect 5160 -3052 5240 -3040
rect 5160 -3108 5172 -3052
rect 5228 -3108 5240 -3052
rect 5160 -3142 5240 -3108
rect 5160 -3198 5172 -3142
rect 5228 -3198 5240 -3142
rect 5160 -3232 5240 -3198
rect 5160 -3288 5172 -3232
rect 5228 -3288 5240 -3232
rect 5160 -3322 5240 -3288
rect 5160 -3378 5172 -3322
rect 5228 -3378 5240 -3322
rect 5160 -3412 5240 -3378
rect 5160 -3468 5172 -3412
rect 5228 -3468 5240 -3412
rect 5160 -3502 5240 -3468
rect 5160 -3558 5172 -3502
rect 5228 -3558 5240 -3502
rect 5160 -3570 5240 -3558
rect 5540 -3052 5620 -3040
rect 5540 -3108 5552 -3052
rect 5608 -3108 5620 -3052
rect 5540 -3142 5620 -3108
rect 5540 -3198 5552 -3142
rect 5608 -3198 5620 -3142
rect 5540 -3232 5620 -3198
rect 5540 -3288 5552 -3232
rect 5608 -3288 5620 -3232
rect 5540 -3322 5620 -3288
rect 5540 -3378 5552 -3322
rect 5608 -3378 5620 -3322
rect 5540 -3412 5620 -3378
rect 5540 -3468 5552 -3412
rect 5608 -3468 5620 -3412
rect 5540 -3502 5620 -3468
rect 5540 -3558 5552 -3502
rect 5608 -3558 5620 -3502
rect 5540 -3570 5620 -3558
rect 5920 -3052 6000 -3040
rect 5920 -3108 5932 -3052
rect 5988 -3108 6000 -3052
rect 5920 -3142 6000 -3108
rect 5920 -3198 5932 -3142
rect 5988 -3198 6000 -3142
rect 5920 -3232 6000 -3198
rect 5920 -3288 5932 -3232
rect 5988 -3288 6000 -3232
rect 5920 -3322 6000 -3288
rect 5920 -3378 5932 -3322
rect 5988 -3378 6000 -3322
rect 5920 -3412 6000 -3378
rect 5920 -3468 5932 -3412
rect 5988 -3468 6000 -3412
rect 5920 -3502 6000 -3468
rect 5920 -3558 5932 -3502
rect 5988 -3558 6000 -3502
rect 5920 -3570 6000 -3558
rect 6300 -3052 6380 -3040
rect 6300 -3108 6312 -3052
rect 6368 -3108 6380 -3052
rect 6300 -3142 6380 -3108
rect 6300 -3198 6312 -3142
rect 6368 -3198 6380 -3142
rect 6300 -3232 6380 -3198
rect 6300 -3288 6312 -3232
rect 6368 -3288 6380 -3232
rect 6300 -3322 6380 -3288
rect 6300 -3378 6312 -3322
rect 6368 -3378 6380 -3322
rect 6300 -3412 6380 -3378
rect 6300 -3468 6312 -3412
rect 6368 -3468 6380 -3412
rect 6300 -3502 6380 -3468
rect 6300 -3558 6312 -3502
rect 6368 -3558 6380 -3502
rect 6300 -3570 6380 -3558
rect 6680 -3052 6760 -3040
rect 6680 -3108 6692 -3052
rect 6748 -3108 6760 -3052
rect 6680 -3142 6760 -3108
rect 6680 -3198 6692 -3142
rect 6748 -3198 6760 -3142
rect 6680 -3232 6760 -3198
rect 6680 -3288 6692 -3232
rect 6748 -3288 6760 -3232
rect 6680 -3322 6760 -3288
rect 6680 -3378 6692 -3322
rect 6748 -3378 6760 -3322
rect 6680 -3412 6760 -3378
rect 6680 -3468 6692 -3412
rect 6748 -3468 6760 -3412
rect 6680 -3502 6760 -3468
rect 6680 -3558 6692 -3502
rect 6748 -3558 6760 -3502
rect 6680 -3570 6760 -3558
rect 7060 -3052 7140 -3040
rect 7060 -3108 7072 -3052
rect 7128 -3108 7140 -3052
rect 7060 -3142 7140 -3108
rect 7060 -3198 7072 -3142
rect 7128 -3198 7140 -3142
rect 7060 -3232 7140 -3198
rect 7060 -3288 7072 -3232
rect 7128 -3288 7140 -3232
rect 7060 -3322 7140 -3288
rect 7060 -3378 7072 -3322
rect 7128 -3378 7140 -3322
rect 7060 -3412 7140 -3378
rect 7060 -3468 7072 -3412
rect 7128 -3468 7140 -3412
rect 7060 -3502 7140 -3468
rect 7060 -3558 7072 -3502
rect 7128 -3558 7140 -3502
rect 7060 -3570 7140 -3558
rect 7440 -3052 7520 -3040
rect 7440 -3108 7452 -3052
rect 7508 -3108 7520 -3052
rect 7440 -3142 7520 -3108
rect 7440 -3198 7452 -3142
rect 7508 -3198 7520 -3142
rect 7440 -3232 7520 -3198
rect 7440 -3288 7452 -3232
rect 7508 -3288 7520 -3232
rect 7440 -3322 7520 -3288
rect 7440 -3378 7452 -3322
rect 7508 -3378 7520 -3322
rect 7440 -3412 7520 -3378
rect 7440 -3468 7452 -3412
rect 7508 -3468 7520 -3412
rect 7440 -3502 7520 -3468
rect 7440 -3558 7452 -3502
rect 7508 -3558 7520 -3502
rect 7440 -3570 7520 -3558
rect 7820 -3052 7900 -3040
rect 7820 -3108 7832 -3052
rect 7888 -3108 7900 -3052
rect 7820 -3142 7900 -3108
rect 7820 -3198 7832 -3142
rect 7888 -3198 7900 -3142
rect 7820 -3232 7900 -3198
rect 7820 -3288 7832 -3232
rect 7888 -3288 7900 -3232
rect 7820 -3322 7900 -3288
rect 7820 -3378 7832 -3322
rect 7888 -3378 7900 -3322
rect 7820 -3412 7900 -3378
rect 7820 -3468 7832 -3412
rect 7888 -3468 7900 -3412
rect 7820 -3502 7900 -3468
rect 7820 -3558 7832 -3502
rect 7888 -3558 7900 -3502
rect 7820 -3570 7900 -3558
rect 8200 -3052 8280 -3040
rect 8200 -3108 8212 -3052
rect 8268 -3108 8280 -3052
rect 8200 -3142 8280 -3108
rect 8200 -3198 8212 -3142
rect 8268 -3198 8280 -3142
rect 8200 -3232 8280 -3198
rect 8200 -3288 8212 -3232
rect 8268 -3288 8280 -3232
rect 8200 -3322 8280 -3288
rect 8200 -3378 8212 -3322
rect 8268 -3378 8280 -3322
rect 8200 -3412 8280 -3378
rect 8200 -3468 8212 -3412
rect 8268 -3468 8280 -3412
rect 8200 -3502 8280 -3468
rect 8200 -3558 8212 -3502
rect 8268 -3558 8280 -3502
rect 8200 -3570 8280 -3558
rect -250 -4214 -170 -4210
rect -250 -4266 -236 -4214
rect -184 -4266 -170 -4214
rect -250 -4290 -170 -4266
rect -250 -4294 2090 -4290
rect -250 -4346 -236 -4294
rect -184 -4346 437 -4294
rect 489 -4346 501 -4294
rect 553 -4346 817 -4294
rect 869 -4346 881 -4294
rect 933 -4346 1197 -4294
rect 1249 -4346 1261 -4294
rect 1313 -4346 1577 -4294
rect 1629 -4346 1641 -4294
rect 1693 -4346 1957 -4294
rect 2009 -4346 2021 -4294
rect 2073 -4346 2090 -4294
rect -250 -4350 2090 -4346
rect 2320 -4294 4190 -4290
rect 2320 -4346 2337 -4294
rect 2389 -4346 2401 -4294
rect 2453 -4346 2717 -4294
rect 2769 -4346 2781 -4294
rect 2833 -4346 3097 -4294
rect 3149 -4346 3161 -4294
rect 3213 -4346 3477 -4294
rect 3529 -4346 3541 -4294
rect 3593 -4346 3857 -4294
rect 3909 -4346 3921 -4294
rect 3973 -4346 4024 -4294
rect 4076 -4302 4124 -4294
rect 4176 -4302 4190 -4294
rect 2320 -4350 4032 -4346
rect 4020 -4358 4032 -4350
rect 4088 -4358 4122 -4302
rect 4178 -4358 4190 -4302
rect 4600 -4294 6470 -4290
rect 4600 -4346 4617 -4294
rect 4669 -4346 4681 -4294
rect 4733 -4346 4997 -4294
rect 5049 -4346 5061 -4294
rect 5113 -4346 5377 -4294
rect 5429 -4346 5441 -4294
rect 5493 -4346 5757 -4294
rect 5809 -4346 5821 -4294
rect 5873 -4346 6137 -4294
rect 6189 -4346 6201 -4294
rect 6253 -4302 6314 -4294
rect 6366 -4302 6404 -4294
rect 6456 -4302 6470 -4294
rect 6253 -4346 6312 -4302
rect 4600 -4350 6312 -4346
rect 4020 -4370 4190 -4358
rect 6300 -4358 6312 -4350
rect 6368 -4358 6402 -4302
rect 6458 -4358 6470 -4302
rect 6500 -4294 8770 -4290
rect 6500 -4346 6517 -4294
rect 6569 -4346 6581 -4294
rect 6633 -4346 6897 -4294
rect 6949 -4346 6961 -4294
rect 7013 -4346 7277 -4294
rect 7329 -4346 7341 -4294
rect 7393 -4346 7657 -4294
rect 7709 -4346 7721 -4294
rect 7773 -4346 8037 -4294
rect 8089 -4346 8101 -4294
rect 8153 -4346 8704 -4294
rect 8756 -4346 8770 -4294
rect 6500 -4350 8770 -4346
rect 6300 -4370 6470 -4358
rect 8690 -4374 8770 -4350
rect 8690 -4426 8704 -4374
rect 8756 -4426 8770 -4374
rect 8690 -4430 8770 -4426
rect 8830 -4662 8910 -4650
rect -250 -4684 -170 -4680
rect -250 -4736 -236 -4684
rect -184 -4736 -170 -4684
rect -250 -4740 -170 -4736
rect 8830 -4718 8842 -4662
rect 8898 -4718 8910 -4662
rect 8830 -4740 8910 -4718
rect -590 -4760 -490 -4750
rect -250 -4752 8910 -4740
rect -590 -4772 -280 -4760
rect -590 -4828 -568 -4772
rect -512 -4828 -280 -4772
rect -250 -4764 8842 -4752
rect -250 -4816 -236 -4764
rect -184 -4808 8842 -4764
rect 8898 -4808 8910 -4752
rect -184 -4816 8910 -4808
rect -250 -4820 8910 -4816
rect -590 -4840 -280 -4828
rect -590 -4850 -490 -4840
rect -360 -4850 -280 -4840
rect -360 -4862 4570 -4850
rect -360 -4918 4032 -4862
rect 4088 -4918 4122 -4862
rect 4178 -4918 4412 -4862
rect 4468 -4918 4502 -4862
rect 4558 -4918 4570 -4862
rect -360 -4930 4570 -4918
rect -590 -4960 -490 -4950
rect -590 -4972 6470 -4960
rect -590 -5028 -568 -4972
rect -512 -5028 232 -4972
rect 288 -5028 322 -4972
rect 378 -5028 6312 -4972
rect 6368 -5028 6402 -4972
rect 6458 -5028 6470 -4972
rect -590 -5040 6470 -5028
rect 8690 -5004 8770 -4990
rect -590 -5050 -490 -5040
rect 8690 -5056 8704 -5004
rect 8756 -5056 8770 -5004
rect 8690 -5070 8770 -5056
rect -350 -5082 8770 -5070
rect -350 -5138 -98 -5082
rect -42 -5138 -8 -5082
rect 48 -5084 8770 -5082
rect 48 -5136 8704 -5084
rect 8756 -5136 8770 -5084
rect 48 -5138 8770 -5136
rect -350 -5150 8770 -5138
rect -590 -5160 -490 -5150
rect -350 -5160 -270 -5150
rect -590 -5172 -270 -5160
rect -590 -5228 -568 -5172
rect -512 -5228 -270 -5172
rect -590 -5240 -270 -5228
rect -590 -5250 -490 -5240
<< via2 >>
rect 4492 5282 4548 5338
rect -238 5032 -182 5088
rect -148 5032 -92 5088
rect 4172 4922 4228 4978
rect 4262 4922 4318 4978
rect 4412 4922 4468 4978
rect 4502 4922 4558 4978
rect -98 4812 -42 4868
rect -8 4812 48 4868
rect 8612 4812 8668 4868
rect 8702 4812 8758 4868
rect 232 4702 288 4758
rect 322 4702 378 4758
rect -98 4242 -42 4298
rect 4172 4262 4228 4318
rect 4262 4262 4318 4318
rect 4522 4316 4578 4318
rect 4522 4264 4524 4316
rect 4524 4264 4576 4316
rect 4576 4264 4578 4316
rect 4522 4262 4578 4264
rect 4612 4311 4668 4318
rect 4612 4262 4614 4311
rect 4614 4262 4666 4311
rect 4666 4262 4668 4311
rect -98 4152 -42 4208
rect 612 3526 668 3528
rect 612 3474 614 3526
rect 614 3474 666 3526
rect 666 3474 668 3526
rect 612 3472 668 3474
rect 612 3436 668 3438
rect 612 3384 614 3436
rect 614 3384 666 3436
rect 666 3384 668 3436
rect 612 3382 668 3384
rect 612 3346 668 3348
rect 612 3294 614 3346
rect 614 3294 666 3346
rect 666 3294 668 3346
rect 612 3292 668 3294
rect 612 3256 668 3258
rect 612 3204 614 3256
rect 614 3204 666 3256
rect 666 3204 668 3256
rect 612 3202 668 3204
rect 612 3166 668 3168
rect 612 3114 614 3166
rect 614 3114 666 3166
rect 666 3114 668 3166
rect 612 3112 668 3114
rect 612 3076 668 3078
rect 612 3024 614 3076
rect 614 3024 666 3076
rect 666 3024 668 3076
rect 612 3022 668 3024
rect 992 3526 1048 3528
rect 992 3474 994 3526
rect 994 3474 1046 3526
rect 1046 3474 1048 3526
rect 992 3472 1048 3474
rect 992 3436 1048 3438
rect 992 3384 994 3436
rect 994 3384 1046 3436
rect 1046 3384 1048 3436
rect 992 3382 1048 3384
rect 992 3346 1048 3348
rect 992 3294 994 3346
rect 994 3294 1046 3346
rect 1046 3294 1048 3346
rect 992 3292 1048 3294
rect 992 3256 1048 3258
rect 992 3204 994 3256
rect 994 3204 1046 3256
rect 1046 3204 1048 3256
rect 992 3202 1048 3204
rect 992 3166 1048 3168
rect 992 3114 994 3166
rect 994 3114 1046 3166
rect 1046 3114 1048 3166
rect 992 3112 1048 3114
rect 992 3076 1048 3078
rect 992 3024 994 3076
rect 994 3024 1046 3076
rect 1046 3024 1048 3076
rect 992 3022 1048 3024
rect 1372 3526 1428 3528
rect 1372 3474 1374 3526
rect 1374 3474 1426 3526
rect 1426 3474 1428 3526
rect 1372 3472 1428 3474
rect 1372 3436 1428 3438
rect 1372 3384 1374 3436
rect 1374 3384 1426 3436
rect 1426 3384 1428 3436
rect 1372 3382 1428 3384
rect 1372 3346 1428 3348
rect 1372 3294 1374 3346
rect 1374 3294 1426 3346
rect 1426 3294 1428 3346
rect 1372 3292 1428 3294
rect 1372 3256 1428 3258
rect 1372 3204 1374 3256
rect 1374 3204 1426 3256
rect 1426 3204 1428 3256
rect 1372 3202 1428 3204
rect 1372 3166 1428 3168
rect 1372 3114 1374 3166
rect 1374 3114 1426 3166
rect 1426 3114 1428 3166
rect 1372 3112 1428 3114
rect 1372 3076 1428 3078
rect 1372 3024 1374 3076
rect 1374 3024 1426 3076
rect 1426 3024 1428 3076
rect 1372 3022 1428 3024
rect 1752 3526 1808 3528
rect 1752 3474 1754 3526
rect 1754 3474 1806 3526
rect 1806 3474 1808 3526
rect 1752 3472 1808 3474
rect 1752 3436 1808 3438
rect 1752 3384 1754 3436
rect 1754 3384 1806 3436
rect 1806 3384 1808 3436
rect 1752 3382 1808 3384
rect 1752 3346 1808 3348
rect 1752 3294 1754 3346
rect 1754 3294 1806 3346
rect 1806 3294 1808 3346
rect 1752 3292 1808 3294
rect 1752 3256 1808 3258
rect 1752 3204 1754 3256
rect 1754 3204 1806 3256
rect 1806 3204 1808 3256
rect 1752 3202 1808 3204
rect 1752 3166 1808 3168
rect 1752 3114 1754 3166
rect 1754 3114 1806 3166
rect 1806 3114 1808 3166
rect 1752 3112 1808 3114
rect 1752 3076 1808 3078
rect 1752 3024 1754 3076
rect 1754 3024 1806 3076
rect 1806 3024 1808 3076
rect 1752 3022 1808 3024
rect 2132 3526 2188 3528
rect 2132 3474 2134 3526
rect 2134 3474 2186 3526
rect 2186 3474 2188 3526
rect 2132 3472 2188 3474
rect 2132 3436 2188 3438
rect 2132 3384 2134 3436
rect 2134 3384 2186 3436
rect 2186 3384 2188 3436
rect 2132 3382 2188 3384
rect 2132 3346 2188 3348
rect 2132 3294 2134 3346
rect 2134 3294 2186 3346
rect 2186 3294 2188 3346
rect 2132 3292 2188 3294
rect 2132 3256 2188 3258
rect 2132 3204 2134 3256
rect 2134 3204 2186 3256
rect 2186 3204 2188 3256
rect 2132 3202 2188 3204
rect 2132 3166 2188 3168
rect 2132 3114 2134 3166
rect 2134 3114 2186 3166
rect 2186 3114 2188 3166
rect 2132 3112 2188 3114
rect 2132 3076 2188 3078
rect 2132 3024 2134 3076
rect 2134 3024 2186 3076
rect 2186 3024 2188 3076
rect 2132 3022 2188 3024
rect 2512 3526 2568 3528
rect 2512 3474 2514 3526
rect 2514 3474 2566 3526
rect 2566 3474 2568 3526
rect 2512 3472 2568 3474
rect 2512 3436 2568 3438
rect 2512 3384 2514 3436
rect 2514 3384 2566 3436
rect 2566 3384 2568 3436
rect 2512 3382 2568 3384
rect 2512 3346 2568 3348
rect 2512 3294 2514 3346
rect 2514 3294 2566 3346
rect 2566 3294 2568 3346
rect 2512 3292 2568 3294
rect 2512 3256 2568 3258
rect 2512 3204 2514 3256
rect 2514 3204 2566 3256
rect 2566 3204 2568 3256
rect 2512 3202 2568 3204
rect 2512 3166 2568 3168
rect 2512 3114 2514 3166
rect 2514 3114 2566 3166
rect 2566 3114 2568 3166
rect 2512 3112 2568 3114
rect 2512 3076 2568 3078
rect 2512 3024 2514 3076
rect 2514 3024 2566 3076
rect 2566 3024 2568 3076
rect 2512 3022 2568 3024
rect 2892 3526 2948 3528
rect 2892 3474 2894 3526
rect 2894 3474 2946 3526
rect 2946 3474 2948 3526
rect 2892 3472 2948 3474
rect 2892 3436 2948 3438
rect 2892 3384 2894 3436
rect 2894 3384 2946 3436
rect 2946 3384 2948 3436
rect 2892 3382 2948 3384
rect 2892 3346 2948 3348
rect 2892 3294 2894 3346
rect 2894 3294 2946 3346
rect 2946 3294 2948 3346
rect 2892 3292 2948 3294
rect 2892 3256 2948 3258
rect 2892 3204 2894 3256
rect 2894 3204 2946 3256
rect 2946 3204 2948 3256
rect 2892 3202 2948 3204
rect 2892 3166 2948 3168
rect 2892 3114 2894 3166
rect 2894 3114 2946 3166
rect 2946 3114 2948 3166
rect 2892 3112 2948 3114
rect 2892 3076 2948 3078
rect 2892 3024 2894 3076
rect 2894 3024 2946 3076
rect 2946 3024 2948 3076
rect 2892 3022 2948 3024
rect 3272 3526 3328 3528
rect 3272 3474 3274 3526
rect 3274 3474 3326 3526
rect 3326 3474 3328 3526
rect 3272 3472 3328 3474
rect 3272 3436 3328 3438
rect 3272 3384 3274 3436
rect 3274 3384 3326 3436
rect 3326 3384 3328 3436
rect 3272 3382 3328 3384
rect 3272 3346 3328 3348
rect 3272 3294 3274 3346
rect 3274 3294 3326 3346
rect 3326 3294 3328 3346
rect 3272 3292 3328 3294
rect 3272 3256 3328 3258
rect 3272 3204 3274 3256
rect 3274 3204 3326 3256
rect 3326 3204 3328 3256
rect 3272 3202 3328 3204
rect 3272 3166 3328 3168
rect 3272 3114 3274 3166
rect 3274 3114 3326 3166
rect 3326 3114 3328 3166
rect 3272 3112 3328 3114
rect 3272 3076 3328 3078
rect 3272 3024 3274 3076
rect 3274 3024 3326 3076
rect 3326 3024 3328 3076
rect 3272 3022 3328 3024
rect 3652 3526 3708 3528
rect 3652 3474 3654 3526
rect 3654 3474 3706 3526
rect 3706 3474 3708 3526
rect 3652 3472 3708 3474
rect 3652 3436 3708 3438
rect 3652 3384 3654 3436
rect 3654 3384 3706 3436
rect 3706 3384 3708 3436
rect 3652 3382 3708 3384
rect 3652 3346 3708 3348
rect 3652 3294 3654 3346
rect 3654 3294 3706 3346
rect 3706 3294 3708 3346
rect 3652 3292 3708 3294
rect 3652 3256 3708 3258
rect 3652 3204 3654 3256
rect 3654 3204 3706 3256
rect 3706 3204 3708 3256
rect 3652 3202 3708 3204
rect 3652 3166 3708 3168
rect 3652 3114 3654 3166
rect 3654 3114 3706 3166
rect 3706 3114 3708 3166
rect 3652 3112 3708 3114
rect 3652 3076 3708 3078
rect 3652 3024 3654 3076
rect 3654 3024 3706 3076
rect 3706 3024 3708 3076
rect 3652 3022 3708 3024
rect 4032 3526 4088 3528
rect 4032 3474 4034 3526
rect 4034 3474 4086 3526
rect 4086 3474 4088 3526
rect 4032 3472 4088 3474
rect 4032 3436 4088 3438
rect 4032 3384 4034 3436
rect 4034 3384 4086 3436
rect 4086 3384 4088 3436
rect 4032 3382 4088 3384
rect 4032 3346 4088 3348
rect 4032 3294 4034 3346
rect 4034 3294 4086 3346
rect 4086 3294 4088 3346
rect 4032 3292 4088 3294
rect 4032 3256 4088 3258
rect 4032 3204 4034 3256
rect 4034 3204 4086 3256
rect 4086 3204 4088 3256
rect 4032 3202 4088 3204
rect 4032 3166 4088 3168
rect 4032 3114 4034 3166
rect 4034 3114 4086 3166
rect 4086 3114 4088 3166
rect 4032 3112 4088 3114
rect 4032 3076 4088 3078
rect 4032 3024 4034 3076
rect 4034 3024 4086 3076
rect 4086 3024 4088 3076
rect 4032 3022 4088 3024
rect -98 2062 -42 2118
rect -98 1972 -42 2028
rect -98 1796 -42 1798
rect -98 1744 -96 1796
rect -96 1744 -44 1796
rect -44 1744 -42 1796
rect -98 1742 -42 1744
rect -98 1706 -42 1708
rect -98 1654 -96 1706
rect -96 1654 -44 1706
rect -44 1654 -42 1706
rect -98 1652 -42 1654
rect 612 1376 668 1378
rect 612 1324 614 1376
rect 614 1324 666 1376
rect 666 1324 668 1376
rect 612 1322 668 1324
rect 612 1286 668 1288
rect 612 1234 614 1286
rect 614 1234 666 1286
rect 666 1234 668 1286
rect 612 1232 668 1234
rect 612 1196 668 1198
rect 612 1144 614 1196
rect 614 1144 666 1196
rect 666 1144 668 1196
rect 612 1142 668 1144
rect 612 1106 668 1108
rect 612 1054 614 1106
rect 614 1054 666 1106
rect 666 1054 668 1106
rect 612 1052 668 1054
rect 612 1016 668 1018
rect 612 964 614 1016
rect 614 964 666 1016
rect 666 964 668 1016
rect 612 962 668 964
rect 612 926 668 928
rect 612 874 614 926
rect 614 874 666 926
rect 666 874 668 926
rect 612 872 668 874
rect 992 1376 1048 1378
rect 992 1324 994 1376
rect 994 1324 1046 1376
rect 1046 1324 1048 1376
rect 992 1322 1048 1324
rect 992 1286 1048 1288
rect 992 1234 994 1286
rect 994 1234 1046 1286
rect 1046 1234 1048 1286
rect 992 1232 1048 1234
rect 992 1196 1048 1198
rect 992 1144 994 1196
rect 994 1144 1046 1196
rect 1046 1144 1048 1196
rect 992 1142 1048 1144
rect 992 1106 1048 1108
rect 992 1054 994 1106
rect 994 1054 1046 1106
rect 1046 1054 1048 1106
rect 992 1052 1048 1054
rect 992 1016 1048 1018
rect 992 964 994 1016
rect 994 964 1046 1016
rect 1046 964 1048 1016
rect 992 962 1048 964
rect 992 926 1048 928
rect 992 874 994 926
rect 994 874 1046 926
rect 1046 874 1048 926
rect 992 872 1048 874
rect 1372 1376 1428 1378
rect 1372 1324 1374 1376
rect 1374 1324 1426 1376
rect 1426 1324 1428 1376
rect 1372 1322 1428 1324
rect 1372 1286 1428 1288
rect 1372 1234 1374 1286
rect 1374 1234 1426 1286
rect 1426 1234 1428 1286
rect 1372 1232 1428 1234
rect 1372 1196 1428 1198
rect 1372 1144 1374 1196
rect 1374 1144 1426 1196
rect 1426 1144 1428 1196
rect 1372 1142 1428 1144
rect 1372 1106 1428 1108
rect 1372 1054 1374 1106
rect 1374 1054 1426 1106
rect 1426 1054 1428 1106
rect 1372 1052 1428 1054
rect 1372 1016 1428 1018
rect 1372 964 1374 1016
rect 1374 964 1426 1016
rect 1426 964 1428 1016
rect 1372 962 1428 964
rect 1372 926 1428 928
rect 1372 874 1374 926
rect 1374 874 1426 926
rect 1426 874 1428 926
rect 1372 872 1428 874
rect 1752 1376 1808 1378
rect 1752 1324 1754 1376
rect 1754 1324 1806 1376
rect 1806 1324 1808 1376
rect 1752 1322 1808 1324
rect 1752 1286 1808 1288
rect 1752 1234 1754 1286
rect 1754 1234 1806 1286
rect 1806 1234 1808 1286
rect 1752 1232 1808 1234
rect 1752 1196 1808 1198
rect 1752 1144 1754 1196
rect 1754 1144 1806 1196
rect 1806 1144 1808 1196
rect 1752 1142 1808 1144
rect 1752 1106 1808 1108
rect 1752 1054 1754 1106
rect 1754 1054 1806 1106
rect 1806 1054 1808 1106
rect 1752 1052 1808 1054
rect 1752 1016 1808 1018
rect 1752 964 1754 1016
rect 1754 964 1806 1016
rect 1806 964 1808 1016
rect 1752 962 1808 964
rect 1752 926 1808 928
rect 1752 874 1754 926
rect 1754 874 1806 926
rect 1806 874 1808 926
rect 1752 872 1808 874
rect 2132 1376 2188 1378
rect 2132 1324 2134 1376
rect 2134 1324 2186 1376
rect 2186 1324 2188 1376
rect 2132 1322 2188 1324
rect 2132 1286 2188 1288
rect 2132 1234 2134 1286
rect 2134 1234 2186 1286
rect 2186 1234 2188 1286
rect 2132 1232 2188 1234
rect 2132 1196 2188 1198
rect 2132 1144 2134 1196
rect 2134 1144 2186 1196
rect 2186 1144 2188 1196
rect 2132 1142 2188 1144
rect 2132 1106 2188 1108
rect 2132 1054 2134 1106
rect 2134 1054 2186 1106
rect 2186 1054 2188 1106
rect 2132 1052 2188 1054
rect 2132 1016 2188 1018
rect 2132 964 2134 1016
rect 2134 964 2186 1016
rect 2186 964 2188 1016
rect 2132 962 2188 964
rect 2132 926 2188 928
rect 2132 874 2134 926
rect 2134 874 2186 926
rect 2186 874 2188 926
rect 2132 872 2188 874
rect 2512 1376 2568 1378
rect 2512 1324 2514 1376
rect 2514 1324 2566 1376
rect 2566 1324 2568 1376
rect 2512 1322 2568 1324
rect 2512 1286 2568 1288
rect 2512 1234 2514 1286
rect 2514 1234 2566 1286
rect 2566 1234 2568 1286
rect 2512 1232 2568 1234
rect 2512 1196 2568 1198
rect 2512 1144 2514 1196
rect 2514 1144 2566 1196
rect 2566 1144 2568 1196
rect 2512 1142 2568 1144
rect 2512 1106 2568 1108
rect 2512 1054 2514 1106
rect 2514 1054 2566 1106
rect 2566 1054 2568 1106
rect 2512 1052 2568 1054
rect 2512 1016 2568 1018
rect 2512 964 2514 1016
rect 2514 964 2566 1016
rect 2566 964 2568 1016
rect 2512 962 2568 964
rect 2512 926 2568 928
rect 2512 874 2514 926
rect 2514 874 2566 926
rect 2566 874 2568 926
rect 2512 872 2568 874
rect 2892 1376 2948 1378
rect 2892 1324 2894 1376
rect 2894 1324 2946 1376
rect 2946 1324 2948 1376
rect 2892 1322 2948 1324
rect 2892 1286 2948 1288
rect 2892 1234 2894 1286
rect 2894 1234 2946 1286
rect 2946 1234 2948 1286
rect 2892 1232 2948 1234
rect 2892 1196 2948 1198
rect 2892 1144 2894 1196
rect 2894 1144 2946 1196
rect 2946 1144 2948 1196
rect 2892 1142 2948 1144
rect 2892 1106 2948 1108
rect 2892 1054 2894 1106
rect 2894 1054 2946 1106
rect 2946 1054 2948 1106
rect 2892 1052 2948 1054
rect 2892 1016 2948 1018
rect 2892 964 2894 1016
rect 2894 964 2946 1016
rect 2946 964 2948 1016
rect 2892 962 2948 964
rect 2892 926 2948 928
rect 2892 874 2894 926
rect 2894 874 2946 926
rect 2946 874 2948 926
rect 2892 872 2948 874
rect 3272 1376 3328 1378
rect 3272 1324 3274 1376
rect 3274 1324 3326 1376
rect 3326 1324 3328 1376
rect 3272 1322 3328 1324
rect 3272 1286 3328 1288
rect 3272 1234 3274 1286
rect 3274 1234 3326 1286
rect 3326 1234 3328 1286
rect 3272 1232 3328 1234
rect 3272 1196 3328 1198
rect 3272 1144 3274 1196
rect 3274 1144 3326 1196
rect 3326 1144 3328 1196
rect 3272 1142 3328 1144
rect 3272 1106 3328 1108
rect 3272 1054 3274 1106
rect 3274 1054 3326 1106
rect 3326 1054 3328 1106
rect 3272 1052 3328 1054
rect 3272 1016 3328 1018
rect 3272 964 3274 1016
rect 3274 964 3326 1016
rect 3326 964 3328 1016
rect 3272 962 3328 964
rect 3272 926 3328 928
rect 3272 874 3274 926
rect 3274 874 3326 926
rect 3326 874 3328 926
rect 3272 872 3328 874
rect 3652 1376 3708 1378
rect 3652 1324 3654 1376
rect 3654 1324 3706 1376
rect 3706 1324 3708 1376
rect 3652 1322 3708 1324
rect 3652 1286 3708 1288
rect 3652 1234 3654 1286
rect 3654 1234 3706 1286
rect 3706 1234 3708 1286
rect 3652 1232 3708 1234
rect 3652 1196 3708 1198
rect 3652 1144 3654 1196
rect 3654 1144 3706 1196
rect 3706 1144 3708 1196
rect 3652 1142 3708 1144
rect 3652 1106 3708 1108
rect 3652 1054 3654 1106
rect 3654 1054 3706 1106
rect 3706 1054 3708 1106
rect 3652 1052 3708 1054
rect 3652 1016 3708 1018
rect 3652 964 3654 1016
rect 3654 964 3706 1016
rect 3706 964 3708 1016
rect 3652 962 3708 964
rect 3652 926 3708 928
rect 3652 874 3654 926
rect 3654 874 3706 926
rect 3706 874 3708 926
rect 3652 872 3708 874
rect 4032 1376 4088 1378
rect 4032 1324 4034 1376
rect 4034 1324 4086 1376
rect 4086 1324 4088 1376
rect 4032 1322 4088 1324
rect 4032 1286 4088 1288
rect 4032 1234 4034 1286
rect 4034 1234 4086 1286
rect 4086 1234 4088 1286
rect 4032 1232 4088 1234
rect 4032 1196 4088 1198
rect 4032 1144 4034 1196
rect 4034 1144 4086 1196
rect 4086 1144 4088 1196
rect 4032 1142 4088 1144
rect 4032 1106 4088 1108
rect 4032 1054 4034 1106
rect 4034 1054 4086 1106
rect 4086 1054 4088 1106
rect 4032 1052 4088 1054
rect 4032 1016 4088 1018
rect 4032 964 4034 1016
rect 4034 964 4086 1016
rect 4086 964 4088 1016
rect 4032 962 4088 964
rect 4032 926 4088 928
rect 4032 874 4034 926
rect 4034 874 4086 926
rect 4086 874 4088 926
rect 4032 872 4088 874
rect -98 112 -42 168
rect -238 -8 -182 48
rect -98 22 -42 78
rect -238 -98 -182 -42
rect 4792 3526 4848 3528
rect 4792 3474 4794 3526
rect 4794 3474 4846 3526
rect 4846 3474 4848 3526
rect 4792 3472 4848 3474
rect 4792 3436 4848 3438
rect 4792 3384 4794 3436
rect 4794 3384 4846 3436
rect 4846 3384 4848 3436
rect 4792 3382 4848 3384
rect 4792 3346 4848 3348
rect 4792 3294 4794 3346
rect 4794 3294 4846 3346
rect 4846 3294 4848 3346
rect 4792 3292 4848 3294
rect 4792 3256 4848 3258
rect 4792 3204 4794 3256
rect 4794 3204 4846 3256
rect 4846 3204 4848 3256
rect 4792 3202 4848 3204
rect 4792 3166 4848 3168
rect 4792 3114 4794 3166
rect 4794 3114 4846 3166
rect 4846 3114 4848 3166
rect 4792 3112 4848 3114
rect 4792 3076 4848 3078
rect 4792 3024 4794 3076
rect 4794 3024 4846 3076
rect 4846 3024 4848 3076
rect 4792 3022 4848 3024
rect 5172 3526 5228 3528
rect 5172 3474 5174 3526
rect 5174 3474 5226 3526
rect 5226 3474 5228 3526
rect 5172 3472 5228 3474
rect 5172 3436 5228 3438
rect 5172 3384 5174 3436
rect 5174 3384 5226 3436
rect 5226 3384 5228 3436
rect 5172 3382 5228 3384
rect 5172 3346 5228 3348
rect 5172 3294 5174 3346
rect 5174 3294 5226 3346
rect 5226 3294 5228 3346
rect 5172 3292 5228 3294
rect 5172 3256 5228 3258
rect 5172 3204 5174 3256
rect 5174 3204 5226 3256
rect 5226 3204 5228 3256
rect 5172 3202 5228 3204
rect 5172 3166 5228 3168
rect 5172 3114 5174 3166
rect 5174 3114 5226 3166
rect 5226 3114 5228 3166
rect 5172 3112 5228 3114
rect 5172 3076 5228 3078
rect 5172 3024 5174 3076
rect 5174 3024 5226 3076
rect 5226 3024 5228 3076
rect 5172 3022 5228 3024
rect 5552 3526 5608 3528
rect 5552 3474 5554 3526
rect 5554 3474 5606 3526
rect 5606 3474 5608 3526
rect 5552 3472 5608 3474
rect 5552 3436 5608 3438
rect 5552 3384 5554 3436
rect 5554 3384 5606 3436
rect 5606 3384 5608 3436
rect 5552 3382 5608 3384
rect 5552 3346 5608 3348
rect 5552 3294 5554 3346
rect 5554 3294 5606 3346
rect 5606 3294 5608 3346
rect 5552 3292 5608 3294
rect 5552 3256 5608 3258
rect 5552 3204 5554 3256
rect 5554 3204 5606 3256
rect 5606 3204 5608 3256
rect 5552 3202 5608 3204
rect 5552 3166 5608 3168
rect 5552 3114 5554 3166
rect 5554 3114 5606 3166
rect 5606 3114 5608 3166
rect 5552 3112 5608 3114
rect 5552 3076 5608 3078
rect 5552 3024 5554 3076
rect 5554 3024 5606 3076
rect 5606 3024 5608 3076
rect 5552 3022 5608 3024
rect 5932 3526 5988 3528
rect 5932 3474 5934 3526
rect 5934 3474 5986 3526
rect 5986 3474 5988 3526
rect 5932 3472 5988 3474
rect 5932 3436 5988 3438
rect 5932 3384 5934 3436
rect 5934 3384 5986 3436
rect 5986 3384 5988 3436
rect 5932 3382 5988 3384
rect 5932 3346 5988 3348
rect 5932 3294 5934 3346
rect 5934 3294 5986 3346
rect 5986 3294 5988 3346
rect 5932 3292 5988 3294
rect 5932 3256 5988 3258
rect 5932 3204 5934 3256
rect 5934 3204 5986 3256
rect 5986 3204 5988 3256
rect 5932 3202 5988 3204
rect 5932 3166 5988 3168
rect 5932 3114 5934 3166
rect 5934 3114 5986 3166
rect 5986 3114 5988 3166
rect 5932 3112 5988 3114
rect 5932 3076 5988 3078
rect 5932 3024 5934 3076
rect 5934 3024 5986 3076
rect 5986 3024 5988 3076
rect 5932 3022 5988 3024
rect 6312 3526 6368 3528
rect 6312 3474 6314 3526
rect 6314 3474 6366 3526
rect 6366 3474 6368 3526
rect 6312 3472 6368 3474
rect 6312 3436 6368 3438
rect 6312 3384 6314 3436
rect 6314 3384 6366 3436
rect 6366 3384 6368 3436
rect 6312 3382 6368 3384
rect 6312 3346 6368 3348
rect 6312 3294 6314 3346
rect 6314 3294 6366 3346
rect 6366 3294 6368 3346
rect 6312 3292 6368 3294
rect 6312 3256 6368 3258
rect 6312 3204 6314 3256
rect 6314 3204 6366 3256
rect 6366 3204 6368 3256
rect 6312 3202 6368 3204
rect 6312 3166 6368 3168
rect 6312 3114 6314 3166
rect 6314 3114 6366 3166
rect 6366 3114 6368 3166
rect 6312 3112 6368 3114
rect 6312 3076 6368 3078
rect 6312 3024 6314 3076
rect 6314 3024 6366 3076
rect 6366 3024 6368 3076
rect 6312 3022 6368 3024
rect 6692 3526 6748 3528
rect 6692 3474 6694 3526
rect 6694 3474 6746 3526
rect 6746 3474 6748 3526
rect 6692 3472 6748 3474
rect 6692 3436 6748 3438
rect 6692 3384 6694 3436
rect 6694 3384 6746 3436
rect 6746 3384 6748 3436
rect 6692 3382 6748 3384
rect 6692 3346 6748 3348
rect 6692 3294 6694 3346
rect 6694 3294 6746 3346
rect 6746 3294 6748 3346
rect 6692 3292 6748 3294
rect 6692 3256 6748 3258
rect 6692 3204 6694 3256
rect 6694 3204 6746 3256
rect 6746 3204 6748 3256
rect 6692 3202 6748 3204
rect 6692 3166 6748 3168
rect 6692 3114 6694 3166
rect 6694 3114 6746 3166
rect 6746 3114 6748 3166
rect 6692 3112 6748 3114
rect 6692 3076 6748 3078
rect 6692 3024 6694 3076
rect 6694 3024 6746 3076
rect 6746 3024 6748 3076
rect 6692 3022 6748 3024
rect 7072 3526 7128 3528
rect 7072 3474 7074 3526
rect 7074 3474 7126 3526
rect 7126 3474 7128 3526
rect 7072 3472 7128 3474
rect 7072 3436 7128 3438
rect 7072 3384 7074 3436
rect 7074 3384 7126 3436
rect 7126 3384 7128 3436
rect 7072 3382 7128 3384
rect 7072 3346 7128 3348
rect 7072 3294 7074 3346
rect 7074 3294 7126 3346
rect 7126 3294 7128 3346
rect 7072 3292 7128 3294
rect 7072 3256 7128 3258
rect 7072 3204 7074 3256
rect 7074 3204 7126 3256
rect 7126 3204 7128 3256
rect 7072 3202 7128 3204
rect 7072 3166 7128 3168
rect 7072 3114 7074 3166
rect 7074 3114 7126 3166
rect 7126 3114 7128 3166
rect 7072 3112 7128 3114
rect 7072 3076 7128 3078
rect 7072 3024 7074 3076
rect 7074 3024 7126 3076
rect 7126 3024 7128 3076
rect 7072 3022 7128 3024
rect 7452 3526 7508 3528
rect 7452 3474 7454 3526
rect 7454 3474 7506 3526
rect 7506 3474 7508 3526
rect 7452 3472 7508 3474
rect 7452 3436 7508 3438
rect 7452 3384 7454 3436
rect 7454 3384 7506 3436
rect 7506 3384 7508 3436
rect 7452 3382 7508 3384
rect 7452 3346 7508 3348
rect 7452 3294 7454 3346
rect 7454 3294 7506 3346
rect 7506 3294 7508 3346
rect 7452 3292 7508 3294
rect 7452 3256 7508 3258
rect 7452 3204 7454 3256
rect 7454 3204 7506 3256
rect 7506 3204 7508 3256
rect 7452 3202 7508 3204
rect 7452 3166 7508 3168
rect 7452 3114 7454 3166
rect 7454 3114 7506 3166
rect 7506 3114 7508 3166
rect 7452 3112 7508 3114
rect 7452 3076 7508 3078
rect 7452 3024 7454 3076
rect 7454 3024 7506 3076
rect 7506 3024 7508 3076
rect 7452 3022 7508 3024
rect 7832 3526 7888 3528
rect 7832 3474 7834 3526
rect 7834 3474 7886 3526
rect 7886 3474 7888 3526
rect 7832 3472 7888 3474
rect 7832 3436 7888 3438
rect 7832 3384 7834 3436
rect 7834 3384 7886 3436
rect 7886 3384 7888 3436
rect 7832 3382 7888 3384
rect 7832 3346 7888 3348
rect 7832 3294 7834 3346
rect 7834 3294 7886 3346
rect 7886 3294 7888 3346
rect 7832 3292 7888 3294
rect 7832 3256 7888 3258
rect 7832 3204 7834 3256
rect 7834 3204 7886 3256
rect 7886 3204 7888 3256
rect 7832 3202 7888 3204
rect 7832 3166 7888 3168
rect 7832 3114 7834 3166
rect 7834 3114 7886 3166
rect 7886 3114 7888 3166
rect 7832 3112 7888 3114
rect 7832 3076 7888 3078
rect 7832 3024 7834 3076
rect 7834 3024 7886 3076
rect 7886 3024 7888 3076
rect 7832 3022 7888 3024
rect 8212 3526 8268 3528
rect 8212 3474 8214 3526
rect 8214 3474 8266 3526
rect 8266 3474 8268 3526
rect 8212 3472 8268 3474
rect 8212 3436 8268 3438
rect 8212 3384 8214 3436
rect 8214 3384 8266 3436
rect 8266 3384 8268 3436
rect 8212 3382 8268 3384
rect 8212 3346 8268 3348
rect 8212 3294 8214 3346
rect 8214 3294 8266 3346
rect 8266 3294 8268 3346
rect 8212 3292 8268 3294
rect 8212 3256 8268 3258
rect 8212 3204 8214 3256
rect 8214 3204 8266 3256
rect 8266 3204 8268 3256
rect 8212 3202 8268 3204
rect 8212 3166 8268 3168
rect 8212 3114 8214 3166
rect 8214 3114 8266 3166
rect 8266 3114 8268 3166
rect 8212 3112 8268 3114
rect 8212 3076 8268 3078
rect 8212 3024 8214 3076
rect 8214 3024 8266 3076
rect 8266 3024 8268 3076
rect 8212 3022 8268 3024
rect 4502 2292 4558 2348
rect 4502 2202 4558 2258
rect 8842 2292 8898 2348
rect 8842 2202 8898 2258
rect 4232 2136 4288 2138
rect 4232 2084 4234 2136
rect 4234 2084 4286 2136
rect 4286 2084 4288 2136
rect 4232 2082 4288 2084
rect 4322 2136 4378 2138
rect 4322 2084 4324 2136
rect 4324 2084 4376 2136
rect 4376 2084 4378 2136
rect 4322 2082 4378 2084
rect 4792 1376 4848 1378
rect 4792 1324 4794 1376
rect 4794 1324 4846 1376
rect 4846 1324 4848 1376
rect 4792 1322 4848 1324
rect 4792 1286 4848 1288
rect 4792 1234 4794 1286
rect 4794 1234 4846 1286
rect 4846 1234 4848 1286
rect 4792 1232 4848 1234
rect 4792 1196 4848 1198
rect 4792 1144 4794 1196
rect 4794 1144 4846 1196
rect 4846 1144 4848 1196
rect 4792 1142 4848 1144
rect 4792 1106 4848 1108
rect 4792 1054 4794 1106
rect 4794 1054 4846 1106
rect 4846 1054 4848 1106
rect 4792 1052 4848 1054
rect 4792 1016 4848 1018
rect 4792 964 4794 1016
rect 4794 964 4846 1016
rect 4846 964 4848 1016
rect 4792 962 4848 964
rect 4792 926 4848 928
rect 4792 874 4794 926
rect 4794 874 4846 926
rect 4846 874 4848 926
rect 4792 872 4848 874
rect 5172 1376 5228 1378
rect 5172 1324 5174 1376
rect 5174 1324 5226 1376
rect 5226 1324 5228 1376
rect 5172 1322 5228 1324
rect 5172 1286 5228 1288
rect 5172 1234 5174 1286
rect 5174 1234 5226 1286
rect 5226 1234 5228 1286
rect 5172 1232 5228 1234
rect 5172 1196 5228 1198
rect 5172 1144 5174 1196
rect 5174 1144 5226 1196
rect 5226 1144 5228 1196
rect 5172 1142 5228 1144
rect 5172 1106 5228 1108
rect 5172 1054 5174 1106
rect 5174 1054 5226 1106
rect 5226 1054 5228 1106
rect 5172 1052 5228 1054
rect 5172 1016 5228 1018
rect 5172 964 5174 1016
rect 5174 964 5226 1016
rect 5226 964 5228 1016
rect 5172 962 5228 964
rect 5172 926 5228 928
rect 5172 874 5174 926
rect 5174 874 5226 926
rect 5226 874 5228 926
rect 5172 872 5228 874
rect 5552 1376 5608 1378
rect 5552 1324 5554 1376
rect 5554 1324 5606 1376
rect 5606 1324 5608 1376
rect 5552 1322 5608 1324
rect 5552 1286 5608 1288
rect 5552 1234 5554 1286
rect 5554 1234 5606 1286
rect 5606 1234 5608 1286
rect 5552 1232 5608 1234
rect 5552 1196 5608 1198
rect 5552 1144 5554 1196
rect 5554 1144 5606 1196
rect 5606 1144 5608 1196
rect 5552 1142 5608 1144
rect 5552 1106 5608 1108
rect 5552 1054 5554 1106
rect 5554 1054 5606 1106
rect 5606 1054 5608 1106
rect 5552 1052 5608 1054
rect 5552 1016 5608 1018
rect 5552 964 5554 1016
rect 5554 964 5606 1016
rect 5606 964 5608 1016
rect 5552 962 5608 964
rect 5552 926 5608 928
rect 5552 874 5554 926
rect 5554 874 5606 926
rect 5606 874 5608 926
rect 5552 872 5608 874
rect 5932 1376 5988 1378
rect 5932 1324 5934 1376
rect 5934 1324 5986 1376
rect 5986 1324 5988 1376
rect 5932 1322 5988 1324
rect 5932 1286 5988 1288
rect 5932 1234 5934 1286
rect 5934 1234 5986 1286
rect 5986 1234 5988 1286
rect 5932 1232 5988 1234
rect 5932 1196 5988 1198
rect 5932 1144 5934 1196
rect 5934 1144 5986 1196
rect 5986 1144 5988 1196
rect 5932 1142 5988 1144
rect 5932 1106 5988 1108
rect 5932 1054 5934 1106
rect 5934 1054 5986 1106
rect 5986 1054 5988 1106
rect 5932 1052 5988 1054
rect 5932 1016 5988 1018
rect 5932 964 5934 1016
rect 5934 964 5986 1016
rect 5986 964 5988 1016
rect 5932 962 5988 964
rect 5932 926 5988 928
rect 5932 874 5934 926
rect 5934 874 5986 926
rect 5986 874 5988 926
rect 5932 872 5988 874
rect 6312 1376 6368 1378
rect 6312 1324 6314 1376
rect 6314 1324 6366 1376
rect 6366 1324 6368 1376
rect 6312 1322 6368 1324
rect 6312 1286 6368 1288
rect 6312 1234 6314 1286
rect 6314 1234 6366 1286
rect 6366 1234 6368 1286
rect 6312 1232 6368 1234
rect 6312 1196 6368 1198
rect 6312 1144 6314 1196
rect 6314 1144 6366 1196
rect 6366 1144 6368 1196
rect 6312 1142 6368 1144
rect 6312 1106 6368 1108
rect 6312 1054 6314 1106
rect 6314 1054 6366 1106
rect 6366 1054 6368 1106
rect 6312 1052 6368 1054
rect 6312 1016 6368 1018
rect 6312 964 6314 1016
rect 6314 964 6366 1016
rect 6366 964 6368 1016
rect 6312 962 6368 964
rect 6312 926 6368 928
rect 6312 874 6314 926
rect 6314 874 6366 926
rect 6366 874 6368 926
rect 6312 872 6368 874
rect 6692 1376 6748 1378
rect 6692 1324 6694 1376
rect 6694 1324 6746 1376
rect 6746 1324 6748 1376
rect 6692 1322 6748 1324
rect 6692 1286 6748 1288
rect 6692 1234 6694 1286
rect 6694 1234 6746 1286
rect 6746 1234 6748 1286
rect 6692 1232 6748 1234
rect 6692 1196 6748 1198
rect 6692 1144 6694 1196
rect 6694 1144 6746 1196
rect 6746 1144 6748 1196
rect 6692 1142 6748 1144
rect 6692 1106 6748 1108
rect 6692 1054 6694 1106
rect 6694 1054 6746 1106
rect 6746 1054 6748 1106
rect 6692 1052 6748 1054
rect 6692 1016 6748 1018
rect 6692 964 6694 1016
rect 6694 964 6746 1016
rect 6746 964 6748 1016
rect 6692 962 6748 964
rect 6692 926 6748 928
rect 6692 874 6694 926
rect 6694 874 6746 926
rect 6746 874 6748 926
rect 6692 872 6748 874
rect 7072 1376 7128 1378
rect 7072 1324 7074 1376
rect 7074 1324 7126 1376
rect 7126 1324 7128 1376
rect 7072 1322 7128 1324
rect 7072 1286 7128 1288
rect 7072 1234 7074 1286
rect 7074 1234 7126 1286
rect 7126 1234 7128 1286
rect 7072 1232 7128 1234
rect 7072 1196 7128 1198
rect 7072 1144 7074 1196
rect 7074 1144 7126 1196
rect 7126 1144 7128 1196
rect 7072 1142 7128 1144
rect 7072 1106 7128 1108
rect 7072 1054 7074 1106
rect 7074 1054 7126 1106
rect 7126 1054 7128 1106
rect 7072 1052 7128 1054
rect 7072 1016 7128 1018
rect 7072 964 7074 1016
rect 7074 964 7126 1016
rect 7126 964 7128 1016
rect 7072 962 7128 964
rect 7072 926 7128 928
rect 7072 874 7074 926
rect 7074 874 7126 926
rect 7126 874 7128 926
rect 7072 872 7128 874
rect 7452 1376 7508 1378
rect 7452 1324 7454 1376
rect 7454 1324 7506 1376
rect 7506 1324 7508 1376
rect 7452 1322 7508 1324
rect 7452 1286 7508 1288
rect 7452 1234 7454 1286
rect 7454 1234 7506 1286
rect 7506 1234 7508 1286
rect 7452 1232 7508 1234
rect 7452 1196 7508 1198
rect 7452 1144 7454 1196
rect 7454 1144 7506 1196
rect 7506 1144 7508 1196
rect 7452 1142 7508 1144
rect 7452 1106 7508 1108
rect 7452 1054 7454 1106
rect 7454 1054 7506 1106
rect 7506 1054 7508 1106
rect 7452 1052 7508 1054
rect 7452 1016 7508 1018
rect 7452 964 7454 1016
rect 7454 964 7506 1016
rect 7506 964 7508 1016
rect 7452 962 7508 964
rect 7452 926 7508 928
rect 7452 874 7454 926
rect 7454 874 7506 926
rect 7506 874 7508 926
rect 7452 872 7508 874
rect 7832 1376 7888 1378
rect 7832 1324 7834 1376
rect 7834 1324 7886 1376
rect 7886 1324 7888 1376
rect 7832 1322 7888 1324
rect 7832 1286 7888 1288
rect 7832 1234 7834 1286
rect 7834 1234 7886 1286
rect 7886 1234 7888 1286
rect 7832 1232 7888 1234
rect 7832 1196 7888 1198
rect 7832 1144 7834 1196
rect 7834 1144 7886 1196
rect 7886 1144 7888 1196
rect 7832 1142 7888 1144
rect 7832 1106 7888 1108
rect 7832 1054 7834 1106
rect 7834 1054 7886 1106
rect 7886 1054 7888 1106
rect 7832 1052 7888 1054
rect 7832 1016 7888 1018
rect 7832 964 7834 1016
rect 7834 964 7886 1016
rect 7886 964 7888 1016
rect 7832 962 7888 964
rect 7832 926 7888 928
rect 7832 874 7834 926
rect 7834 874 7886 926
rect 7886 874 7888 926
rect 7832 872 7888 874
rect 8212 1376 8268 1378
rect 8212 1324 8214 1376
rect 8214 1324 8266 1376
rect 8266 1324 8268 1376
rect 8212 1322 8268 1324
rect 8212 1286 8268 1288
rect 8212 1234 8214 1286
rect 8214 1234 8266 1286
rect 8266 1234 8268 1286
rect 8212 1232 8268 1234
rect 8212 1196 8268 1198
rect 8212 1144 8214 1196
rect 8214 1144 8266 1196
rect 8266 1144 8268 1196
rect 8212 1142 8268 1144
rect 8212 1106 8268 1108
rect 8212 1054 8214 1106
rect 8214 1054 8266 1106
rect 8266 1054 8268 1106
rect 8212 1052 8268 1054
rect 8212 1016 8268 1018
rect 8212 964 8214 1016
rect 8214 964 8266 1016
rect 8266 964 8268 1016
rect 8212 962 8268 964
rect 8212 926 8268 928
rect 8212 874 8214 926
rect 8214 874 8266 926
rect 8266 874 8268 926
rect 8212 872 8268 874
rect 4502 112 4558 168
rect 4502 22 4558 78
rect 8842 112 8898 168
rect 8842 22 8898 78
rect 612 -864 668 -862
rect 612 -916 614 -864
rect 614 -916 666 -864
rect 666 -916 668 -864
rect 612 -918 668 -916
rect 612 -954 668 -952
rect 612 -1006 614 -954
rect 614 -1006 666 -954
rect 666 -1006 668 -954
rect 612 -1008 668 -1006
rect 612 -1044 668 -1042
rect 612 -1096 614 -1044
rect 614 -1096 666 -1044
rect 666 -1096 668 -1044
rect 612 -1098 668 -1096
rect 612 -1134 668 -1132
rect 612 -1186 614 -1134
rect 614 -1186 666 -1134
rect 666 -1186 668 -1134
rect 612 -1188 668 -1186
rect 612 -1224 668 -1222
rect 612 -1276 614 -1224
rect 614 -1276 666 -1224
rect 666 -1276 668 -1224
rect 612 -1278 668 -1276
rect 612 -1314 668 -1312
rect 612 -1366 614 -1314
rect 614 -1366 666 -1314
rect 666 -1366 668 -1314
rect 612 -1368 668 -1366
rect 992 -864 1048 -862
rect 992 -916 994 -864
rect 994 -916 1046 -864
rect 1046 -916 1048 -864
rect 992 -918 1048 -916
rect 992 -954 1048 -952
rect 992 -1006 994 -954
rect 994 -1006 1046 -954
rect 1046 -1006 1048 -954
rect 992 -1008 1048 -1006
rect 992 -1044 1048 -1042
rect 992 -1096 994 -1044
rect 994 -1096 1046 -1044
rect 1046 -1096 1048 -1044
rect 992 -1098 1048 -1096
rect 992 -1134 1048 -1132
rect 992 -1186 994 -1134
rect 994 -1186 1046 -1134
rect 1046 -1186 1048 -1134
rect 992 -1188 1048 -1186
rect 992 -1224 1048 -1222
rect 992 -1276 994 -1224
rect 994 -1276 1046 -1224
rect 1046 -1276 1048 -1224
rect 992 -1278 1048 -1276
rect 992 -1314 1048 -1312
rect 992 -1366 994 -1314
rect 994 -1366 1046 -1314
rect 1046 -1366 1048 -1314
rect 992 -1368 1048 -1366
rect 1372 -864 1428 -862
rect 1372 -916 1374 -864
rect 1374 -916 1426 -864
rect 1426 -916 1428 -864
rect 1372 -918 1428 -916
rect 1372 -954 1428 -952
rect 1372 -1006 1374 -954
rect 1374 -1006 1426 -954
rect 1426 -1006 1428 -954
rect 1372 -1008 1428 -1006
rect 1372 -1044 1428 -1042
rect 1372 -1096 1374 -1044
rect 1374 -1096 1426 -1044
rect 1426 -1096 1428 -1044
rect 1372 -1098 1428 -1096
rect 1372 -1134 1428 -1132
rect 1372 -1186 1374 -1134
rect 1374 -1186 1426 -1134
rect 1426 -1186 1428 -1134
rect 1372 -1188 1428 -1186
rect 1372 -1224 1428 -1222
rect 1372 -1276 1374 -1224
rect 1374 -1276 1426 -1224
rect 1426 -1276 1428 -1224
rect 1372 -1278 1428 -1276
rect 1372 -1314 1428 -1312
rect 1372 -1366 1374 -1314
rect 1374 -1366 1426 -1314
rect 1426 -1366 1428 -1314
rect 1372 -1368 1428 -1366
rect 1752 -864 1808 -862
rect 1752 -916 1754 -864
rect 1754 -916 1806 -864
rect 1806 -916 1808 -864
rect 1752 -918 1808 -916
rect 1752 -954 1808 -952
rect 1752 -1006 1754 -954
rect 1754 -1006 1806 -954
rect 1806 -1006 1808 -954
rect 1752 -1008 1808 -1006
rect 1752 -1044 1808 -1042
rect 1752 -1096 1754 -1044
rect 1754 -1096 1806 -1044
rect 1806 -1096 1808 -1044
rect 1752 -1098 1808 -1096
rect 1752 -1134 1808 -1132
rect 1752 -1186 1754 -1134
rect 1754 -1186 1806 -1134
rect 1806 -1186 1808 -1134
rect 1752 -1188 1808 -1186
rect 1752 -1224 1808 -1222
rect 1752 -1276 1754 -1224
rect 1754 -1276 1806 -1224
rect 1806 -1276 1808 -1224
rect 1752 -1278 1808 -1276
rect 1752 -1314 1808 -1312
rect 1752 -1366 1754 -1314
rect 1754 -1366 1806 -1314
rect 1806 -1366 1808 -1314
rect 1752 -1368 1808 -1366
rect 2132 -864 2188 -862
rect 2132 -916 2134 -864
rect 2134 -916 2186 -864
rect 2186 -916 2188 -864
rect 2132 -918 2188 -916
rect 2132 -954 2188 -952
rect 2132 -1006 2134 -954
rect 2134 -1006 2186 -954
rect 2186 -1006 2188 -954
rect 2132 -1008 2188 -1006
rect 2132 -1044 2188 -1042
rect 2132 -1096 2134 -1044
rect 2134 -1096 2186 -1044
rect 2186 -1096 2188 -1044
rect 2132 -1098 2188 -1096
rect 2132 -1134 2188 -1132
rect 2132 -1186 2134 -1134
rect 2134 -1186 2186 -1134
rect 2186 -1186 2188 -1134
rect 2132 -1188 2188 -1186
rect 2132 -1224 2188 -1222
rect 2132 -1276 2134 -1224
rect 2134 -1276 2186 -1224
rect 2186 -1276 2188 -1224
rect 2132 -1278 2188 -1276
rect 2132 -1314 2188 -1312
rect 2132 -1366 2134 -1314
rect 2134 -1366 2186 -1314
rect 2186 -1366 2188 -1314
rect 2132 -1368 2188 -1366
rect 2512 -864 2568 -862
rect 2512 -916 2514 -864
rect 2514 -916 2566 -864
rect 2566 -916 2568 -864
rect 2512 -918 2568 -916
rect 2512 -954 2568 -952
rect 2512 -1006 2514 -954
rect 2514 -1006 2566 -954
rect 2566 -1006 2568 -954
rect 2512 -1008 2568 -1006
rect 2512 -1044 2568 -1042
rect 2512 -1096 2514 -1044
rect 2514 -1096 2566 -1044
rect 2566 -1096 2568 -1044
rect 2512 -1098 2568 -1096
rect 2512 -1134 2568 -1132
rect 2512 -1186 2514 -1134
rect 2514 -1186 2566 -1134
rect 2566 -1186 2568 -1134
rect 2512 -1188 2568 -1186
rect 2512 -1224 2568 -1222
rect 2512 -1276 2514 -1224
rect 2514 -1276 2566 -1224
rect 2566 -1276 2568 -1224
rect 2512 -1278 2568 -1276
rect 2512 -1314 2568 -1312
rect 2512 -1366 2514 -1314
rect 2514 -1366 2566 -1314
rect 2566 -1366 2568 -1314
rect 2512 -1368 2568 -1366
rect 2892 -864 2948 -862
rect 2892 -916 2894 -864
rect 2894 -916 2946 -864
rect 2946 -916 2948 -864
rect 2892 -918 2948 -916
rect 2892 -954 2948 -952
rect 2892 -1006 2894 -954
rect 2894 -1006 2946 -954
rect 2946 -1006 2948 -954
rect 2892 -1008 2948 -1006
rect 2892 -1044 2948 -1042
rect 2892 -1096 2894 -1044
rect 2894 -1096 2946 -1044
rect 2946 -1096 2948 -1044
rect 2892 -1098 2948 -1096
rect 2892 -1134 2948 -1132
rect 2892 -1186 2894 -1134
rect 2894 -1186 2946 -1134
rect 2946 -1186 2948 -1134
rect 2892 -1188 2948 -1186
rect 2892 -1224 2948 -1222
rect 2892 -1276 2894 -1224
rect 2894 -1276 2946 -1224
rect 2946 -1276 2948 -1224
rect 2892 -1278 2948 -1276
rect 2892 -1314 2948 -1312
rect 2892 -1366 2894 -1314
rect 2894 -1366 2946 -1314
rect 2946 -1366 2948 -1314
rect 2892 -1368 2948 -1366
rect 3272 -864 3328 -862
rect 3272 -916 3274 -864
rect 3274 -916 3326 -864
rect 3326 -916 3328 -864
rect 3272 -918 3328 -916
rect 3272 -954 3328 -952
rect 3272 -1006 3274 -954
rect 3274 -1006 3326 -954
rect 3326 -1006 3328 -954
rect 3272 -1008 3328 -1006
rect 3272 -1044 3328 -1042
rect 3272 -1096 3274 -1044
rect 3274 -1096 3326 -1044
rect 3326 -1096 3328 -1044
rect 3272 -1098 3328 -1096
rect 3272 -1134 3328 -1132
rect 3272 -1186 3274 -1134
rect 3274 -1186 3326 -1134
rect 3326 -1186 3328 -1134
rect 3272 -1188 3328 -1186
rect 3272 -1224 3328 -1222
rect 3272 -1276 3274 -1224
rect 3274 -1276 3326 -1224
rect 3326 -1276 3328 -1224
rect 3272 -1278 3328 -1276
rect 3272 -1314 3328 -1312
rect 3272 -1366 3274 -1314
rect 3274 -1366 3326 -1314
rect 3326 -1366 3328 -1314
rect 3272 -1368 3328 -1366
rect 3652 -864 3708 -862
rect 3652 -916 3654 -864
rect 3654 -916 3706 -864
rect 3706 -916 3708 -864
rect 3652 -918 3708 -916
rect 3652 -954 3708 -952
rect 3652 -1006 3654 -954
rect 3654 -1006 3706 -954
rect 3706 -1006 3708 -954
rect 3652 -1008 3708 -1006
rect 3652 -1044 3708 -1042
rect 3652 -1096 3654 -1044
rect 3654 -1096 3706 -1044
rect 3706 -1096 3708 -1044
rect 3652 -1098 3708 -1096
rect 3652 -1134 3708 -1132
rect 3652 -1186 3654 -1134
rect 3654 -1186 3706 -1134
rect 3706 -1186 3708 -1134
rect 3652 -1188 3708 -1186
rect 3652 -1224 3708 -1222
rect 3652 -1276 3654 -1224
rect 3654 -1276 3706 -1224
rect 3706 -1276 3708 -1224
rect 3652 -1278 3708 -1276
rect 3652 -1314 3708 -1312
rect 3652 -1366 3654 -1314
rect 3654 -1366 3706 -1314
rect 3706 -1366 3708 -1314
rect 3652 -1368 3708 -1366
rect 4032 -864 4088 -862
rect 4032 -916 4034 -864
rect 4034 -916 4086 -864
rect 4086 -916 4088 -864
rect 4032 -918 4088 -916
rect 4032 -954 4088 -952
rect 4032 -1006 4034 -954
rect 4034 -1006 4086 -954
rect 4086 -1006 4088 -954
rect 4032 -1008 4088 -1006
rect 4032 -1044 4088 -1042
rect 4032 -1096 4034 -1044
rect 4034 -1096 4086 -1044
rect 4086 -1096 4088 -1044
rect 4032 -1098 4088 -1096
rect 4032 -1134 4088 -1132
rect 4032 -1186 4034 -1134
rect 4034 -1186 4086 -1134
rect 4086 -1186 4088 -1134
rect 4032 -1188 4088 -1186
rect 4032 -1224 4088 -1222
rect 4032 -1276 4034 -1224
rect 4034 -1276 4086 -1224
rect 4086 -1276 4088 -1224
rect 4032 -1278 4088 -1276
rect 4032 -1314 4088 -1312
rect 4032 -1366 4034 -1314
rect 4034 -1366 4086 -1314
rect 4086 -1366 4088 -1314
rect 4032 -1368 4088 -1366
rect -568 -2168 -512 -2112
rect 8702 -118 8758 -62
rect 8702 -208 8758 -152
rect 4792 -864 4848 -862
rect 4792 -916 4794 -864
rect 4794 -916 4846 -864
rect 4846 -916 4848 -864
rect 4792 -918 4848 -916
rect 4792 -954 4848 -952
rect 4792 -1006 4794 -954
rect 4794 -1006 4846 -954
rect 4846 -1006 4848 -954
rect 4792 -1008 4848 -1006
rect 4792 -1044 4848 -1042
rect 4792 -1096 4794 -1044
rect 4794 -1096 4846 -1044
rect 4846 -1096 4848 -1044
rect 4792 -1098 4848 -1096
rect 4792 -1134 4848 -1132
rect 4792 -1186 4794 -1134
rect 4794 -1186 4846 -1134
rect 4846 -1186 4848 -1134
rect 4792 -1188 4848 -1186
rect 4792 -1224 4848 -1222
rect 4792 -1276 4794 -1224
rect 4794 -1276 4846 -1224
rect 4846 -1276 4848 -1224
rect 4792 -1278 4848 -1276
rect 4792 -1314 4848 -1312
rect 4792 -1366 4794 -1314
rect 4794 -1366 4846 -1314
rect 4846 -1366 4848 -1314
rect 4792 -1368 4848 -1366
rect 5172 -864 5228 -862
rect 5172 -916 5174 -864
rect 5174 -916 5226 -864
rect 5226 -916 5228 -864
rect 5172 -918 5228 -916
rect 5172 -954 5228 -952
rect 5172 -1006 5174 -954
rect 5174 -1006 5226 -954
rect 5226 -1006 5228 -954
rect 5172 -1008 5228 -1006
rect 5172 -1044 5228 -1042
rect 5172 -1096 5174 -1044
rect 5174 -1096 5226 -1044
rect 5226 -1096 5228 -1044
rect 5172 -1098 5228 -1096
rect 5172 -1134 5228 -1132
rect 5172 -1186 5174 -1134
rect 5174 -1186 5226 -1134
rect 5226 -1186 5228 -1134
rect 5172 -1188 5228 -1186
rect 5172 -1224 5228 -1222
rect 5172 -1276 5174 -1224
rect 5174 -1276 5226 -1224
rect 5226 -1276 5228 -1224
rect 5172 -1278 5228 -1276
rect 5172 -1314 5228 -1312
rect 5172 -1366 5174 -1314
rect 5174 -1366 5226 -1314
rect 5226 -1366 5228 -1314
rect 5172 -1368 5228 -1366
rect 5552 -864 5608 -862
rect 5552 -916 5554 -864
rect 5554 -916 5606 -864
rect 5606 -916 5608 -864
rect 5552 -918 5608 -916
rect 5552 -954 5608 -952
rect 5552 -1006 5554 -954
rect 5554 -1006 5606 -954
rect 5606 -1006 5608 -954
rect 5552 -1008 5608 -1006
rect 5552 -1044 5608 -1042
rect 5552 -1096 5554 -1044
rect 5554 -1096 5606 -1044
rect 5606 -1096 5608 -1044
rect 5552 -1098 5608 -1096
rect 5552 -1134 5608 -1132
rect 5552 -1186 5554 -1134
rect 5554 -1186 5606 -1134
rect 5606 -1186 5608 -1134
rect 5552 -1188 5608 -1186
rect 5552 -1224 5608 -1222
rect 5552 -1276 5554 -1224
rect 5554 -1276 5606 -1224
rect 5606 -1276 5608 -1224
rect 5552 -1278 5608 -1276
rect 5552 -1314 5608 -1312
rect 5552 -1366 5554 -1314
rect 5554 -1366 5606 -1314
rect 5606 -1366 5608 -1314
rect 5552 -1368 5608 -1366
rect 5932 -864 5988 -862
rect 5932 -916 5934 -864
rect 5934 -916 5986 -864
rect 5986 -916 5988 -864
rect 5932 -918 5988 -916
rect 5932 -954 5988 -952
rect 5932 -1006 5934 -954
rect 5934 -1006 5986 -954
rect 5986 -1006 5988 -954
rect 5932 -1008 5988 -1006
rect 5932 -1044 5988 -1042
rect 5932 -1096 5934 -1044
rect 5934 -1096 5986 -1044
rect 5986 -1096 5988 -1044
rect 5932 -1098 5988 -1096
rect 5932 -1134 5988 -1132
rect 5932 -1186 5934 -1134
rect 5934 -1186 5986 -1134
rect 5986 -1186 5988 -1134
rect 5932 -1188 5988 -1186
rect 5932 -1224 5988 -1222
rect 5932 -1276 5934 -1224
rect 5934 -1276 5986 -1224
rect 5986 -1276 5988 -1224
rect 5932 -1278 5988 -1276
rect 5932 -1314 5988 -1312
rect 5932 -1366 5934 -1314
rect 5934 -1366 5986 -1314
rect 5986 -1366 5988 -1314
rect 5932 -1368 5988 -1366
rect 6312 -864 6368 -862
rect 6312 -916 6314 -864
rect 6314 -916 6366 -864
rect 6366 -916 6368 -864
rect 6312 -918 6368 -916
rect 6312 -954 6368 -952
rect 6312 -1006 6314 -954
rect 6314 -1006 6366 -954
rect 6366 -1006 6368 -954
rect 6312 -1008 6368 -1006
rect 6312 -1044 6368 -1042
rect 6312 -1096 6314 -1044
rect 6314 -1096 6366 -1044
rect 6366 -1096 6368 -1044
rect 6312 -1098 6368 -1096
rect 6312 -1134 6368 -1132
rect 6312 -1186 6314 -1134
rect 6314 -1186 6366 -1134
rect 6366 -1186 6368 -1134
rect 6312 -1188 6368 -1186
rect 6312 -1224 6368 -1222
rect 6312 -1276 6314 -1224
rect 6314 -1276 6366 -1224
rect 6366 -1276 6368 -1224
rect 6312 -1278 6368 -1276
rect 6312 -1314 6368 -1312
rect 6312 -1366 6314 -1314
rect 6314 -1366 6366 -1314
rect 6366 -1366 6368 -1314
rect 6312 -1368 6368 -1366
rect 6692 -864 6748 -862
rect 6692 -916 6694 -864
rect 6694 -916 6746 -864
rect 6746 -916 6748 -864
rect 6692 -918 6748 -916
rect 6692 -954 6748 -952
rect 6692 -1006 6694 -954
rect 6694 -1006 6746 -954
rect 6746 -1006 6748 -954
rect 6692 -1008 6748 -1006
rect 6692 -1044 6748 -1042
rect 6692 -1096 6694 -1044
rect 6694 -1096 6746 -1044
rect 6746 -1096 6748 -1044
rect 6692 -1098 6748 -1096
rect 6692 -1134 6748 -1132
rect 6692 -1186 6694 -1134
rect 6694 -1186 6746 -1134
rect 6746 -1186 6748 -1134
rect 6692 -1188 6748 -1186
rect 6692 -1224 6748 -1222
rect 6692 -1276 6694 -1224
rect 6694 -1276 6746 -1224
rect 6746 -1276 6748 -1224
rect 6692 -1278 6748 -1276
rect 6692 -1314 6748 -1312
rect 6692 -1366 6694 -1314
rect 6694 -1366 6746 -1314
rect 6746 -1366 6748 -1314
rect 6692 -1368 6748 -1366
rect 7072 -864 7128 -862
rect 7072 -916 7074 -864
rect 7074 -916 7126 -864
rect 7126 -916 7128 -864
rect 7072 -918 7128 -916
rect 7072 -954 7128 -952
rect 7072 -1006 7074 -954
rect 7074 -1006 7126 -954
rect 7126 -1006 7128 -954
rect 7072 -1008 7128 -1006
rect 7072 -1044 7128 -1042
rect 7072 -1096 7074 -1044
rect 7074 -1096 7126 -1044
rect 7126 -1096 7128 -1044
rect 7072 -1098 7128 -1096
rect 7072 -1134 7128 -1132
rect 7072 -1186 7074 -1134
rect 7074 -1186 7126 -1134
rect 7126 -1186 7128 -1134
rect 7072 -1188 7128 -1186
rect 7072 -1224 7128 -1222
rect 7072 -1276 7074 -1224
rect 7074 -1276 7126 -1224
rect 7126 -1276 7128 -1224
rect 7072 -1278 7128 -1276
rect 7072 -1314 7128 -1312
rect 7072 -1366 7074 -1314
rect 7074 -1366 7126 -1314
rect 7126 -1366 7128 -1314
rect 7072 -1368 7128 -1366
rect 7452 -864 7508 -862
rect 7452 -916 7454 -864
rect 7454 -916 7506 -864
rect 7506 -916 7508 -864
rect 7452 -918 7508 -916
rect 7452 -954 7508 -952
rect 7452 -1006 7454 -954
rect 7454 -1006 7506 -954
rect 7506 -1006 7508 -954
rect 7452 -1008 7508 -1006
rect 7452 -1044 7508 -1042
rect 7452 -1096 7454 -1044
rect 7454 -1096 7506 -1044
rect 7506 -1096 7508 -1044
rect 7452 -1098 7508 -1096
rect 7452 -1134 7508 -1132
rect 7452 -1186 7454 -1134
rect 7454 -1186 7506 -1134
rect 7506 -1186 7508 -1134
rect 7452 -1188 7508 -1186
rect 7452 -1224 7508 -1222
rect 7452 -1276 7454 -1224
rect 7454 -1276 7506 -1224
rect 7506 -1276 7508 -1224
rect 7452 -1278 7508 -1276
rect 7452 -1314 7508 -1312
rect 7452 -1366 7454 -1314
rect 7454 -1366 7506 -1314
rect 7506 -1366 7508 -1314
rect 7452 -1368 7508 -1366
rect 7832 -864 7888 -862
rect 7832 -916 7834 -864
rect 7834 -916 7886 -864
rect 7886 -916 7888 -864
rect 7832 -918 7888 -916
rect 7832 -954 7888 -952
rect 7832 -1006 7834 -954
rect 7834 -1006 7886 -954
rect 7886 -1006 7888 -954
rect 7832 -1008 7888 -1006
rect 7832 -1044 7888 -1042
rect 7832 -1096 7834 -1044
rect 7834 -1096 7886 -1044
rect 7886 -1096 7888 -1044
rect 7832 -1098 7888 -1096
rect 7832 -1134 7888 -1132
rect 7832 -1186 7834 -1134
rect 7834 -1186 7886 -1134
rect 7886 -1186 7888 -1134
rect 7832 -1188 7888 -1186
rect 7832 -1224 7888 -1222
rect 7832 -1276 7834 -1224
rect 7834 -1276 7886 -1224
rect 7886 -1276 7888 -1224
rect 7832 -1278 7888 -1276
rect 7832 -1314 7888 -1312
rect 7832 -1366 7834 -1314
rect 7834 -1366 7886 -1314
rect 7886 -1366 7888 -1314
rect 7832 -1368 7888 -1366
rect 8212 -864 8268 -862
rect 8212 -916 8214 -864
rect 8214 -916 8266 -864
rect 8266 -916 8268 -864
rect 8212 -918 8268 -916
rect 8212 -954 8268 -952
rect 8212 -1006 8214 -954
rect 8214 -1006 8266 -954
rect 8266 -1006 8268 -954
rect 8212 -1008 8268 -1006
rect 8212 -1044 8268 -1042
rect 8212 -1096 8214 -1044
rect 8214 -1096 8266 -1044
rect 8266 -1096 8268 -1044
rect 8212 -1098 8268 -1096
rect 8212 -1134 8268 -1132
rect 8212 -1186 8214 -1134
rect 8214 -1186 8266 -1134
rect 8266 -1186 8268 -1134
rect 8212 -1188 8268 -1186
rect 8212 -1224 8268 -1222
rect 8212 -1276 8214 -1224
rect 8214 -1276 8266 -1224
rect 8266 -1276 8268 -1224
rect 8212 -1278 8268 -1276
rect 8212 -1314 8268 -1312
rect 8212 -1366 8214 -1314
rect 8214 -1366 8266 -1314
rect 8266 -1366 8268 -1314
rect 8212 -1368 8268 -1366
rect -238 -2298 -182 -2242
rect -238 -2388 -182 -2332
rect 8702 -2298 8758 -2242
rect 8702 -2388 8758 -2332
rect 612 -3054 668 -3052
rect 612 -3106 614 -3054
rect 614 -3106 666 -3054
rect 666 -3106 668 -3054
rect 612 -3108 668 -3106
rect 612 -3144 668 -3142
rect 612 -3196 614 -3144
rect 614 -3196 666 -3144
rect 666 -3196 668 -3144
rect 612 -3198 668 -3196
rect 612 -3234 668 -3232
rect 612 -3286 614 -3234
rect 614 -3286 666 -3234
rect 666 -3286 668 -3234
rect 612 -3288 668 -3286
rect 612 -3324 668 -3322
rect 612 -3376 614 -3324
rect 614 -3376 666 -3324
rect 666 -3376 668 -3324
rect 612 -3378 668 -3376
rect 612 -3414 668 -3412
rect 612 -3466 614 -3414
rect 614 -3466 666 -3414
rect 666 -3466 668 -3414
rect 612 -3468 668 -3466
rect 612 -3504 668 -3502
rect 612 -3556 614 -3504
rect 614 -3556 666 -3504
rect 666 -3556 668 -3504
rect 612 -3558 668 -3556
rect 992 -3054 1048 -3052
rect 992 -3106 994 -3054
rect 994 -3106 1046 -3054
rect 1046 -3106 1048 -3054
rect 992 -3108 1048 -3106
rect 992 -3144 1048 -3142
rect 992 -3196 994 -3144
rect 994 -3196 1046 -3144
rect 1046 -3196 1048 -3144
rect 992 -3198 1048 -3196
rect 992 -3234 1048 -3232
rect 992 -3286 994 -3234
rect 994 -3286 1046 -3234
rect 1046 -3286 1048 -3234
rect 992 -3288 1048 -3286
rect 992 -3324 1048 -3322
rect 992 -3376 994 -3324
rect 994 -3376 1046 -3324
rect 1046 -3376 1048 -3324
rect 992 -3378 1048 -3376
rect 992 -3414 1048 -3412
rect 992 -3466 994 -3414
rect 994 -3466 1046 -3414
rect 1046 -3466 1048 -3414
rect 992 -3468 1048 -3466
rect 992 -3504 1048 -3502
rect 992 -3556 994 -3504
rect 994 -3556 1046 -3504
rect 1046 -3556 1048 -3504
rect 992 -3558 1048 -3556
rect 1372 -3054 1428 -3052
rect 1372 -3106 1374 -3054
rect 1374 -3106 1426 -3054
rect 1426 -3106 1428 -3054
rect 1372 -3108 1428 -3106
rect 1372 -3144 1428 -3142
rect 1372 -3196 1374 -3144
rect 1374 -3196 1426 -3144
rect 1426 -3196 1428 -3144
rect 1372 -3198 1428 -3196
rect 1372 -3234 1428 -3232
rect 1372 -3286 1374 -3234
rect 1374 -3286 1426 -3234
rect 1426 -3286 1428 -3234
rect 1372 -3288 1428 -3286
rect 1372 -3324 1428 -3322
rect 1372 -3376 1374 -3324
rect 1374 -3376 1426 -3324
rect 1426 -3376 1428 -3324
rect 1372 -3378 1428 -3376
rect 1372 -3414 1428 -3412
rect 1372 -3466 1374 -3414
rect 1374 -3466 1426 -3414
rect 1426 -3466 1428 -3414
rect 1372 -3468 1428 -3466
rect 1372 -3504 1428 -3502
rect 1372 -3556 1374 -3504
rect 1374 -3556 1426 -3504
rect 1426 -3556 1428 -3504
rect 1372 -3558 1428 -3556
rect 1752 -3054 1808 -3052
rect 1752 -3106 1754 -3054
rect 1754 -3106 1806 -3054
rect 1806 -3106 1808 -3054
rect 1752 -3108 1808 -3106
rect 1752 -3144 1808 -3142
rect 1752 -3196 1754 -3144
rect 1754 -3196 1806 -3144
rect 1806 -3196 1808 -3144
rect 1752 -3198 1808 -3196
rect 1752 -3234 1808 -3232
rect 1752 -3286 1754 -3234
rect 1754 -3286 1806 -3234
rect 1806 -3286 1808 -3234
rect 1752 -3288 1808 -3286
rect 1752 -3324 1808 -3322
rect 1752 -3376 1754 -3324
rect 1754 -3376 1806 -3324
rect 1806 -3376 1808 -3324
rect 1752 -3378 1808 -3376
rect 1752 -3414 1808 -3412
rect 1752 -3466 1754 -3414
rect 1754 -3466 1806 -3414
rect 1806 -3466 1808 -3414
rect 1752 -3468 1808 -3466
rect 1752 -3504 1808 -3502
rect 1752 -3556 1754 -3504
rect 1754 -3556 1806 -3504
rect 1806 -3556 1808 -3504
rect 1752 -3558 1808 -3556
rect 2132 -3054 2188 -3052
rect 2132 -3106 2134 -3054
rect 2134 -3106 2186 -3054
rect 2186 -3106 2188 -3054
rect 2132 -3108 2188 -3106
rect 2132 -3144 2188 -3142
rect 2132 -3196 2134 -3144
rect 2134 -3196 2186 -3144
rect 2186 -3196 2188 -3144
rect 2132 -3198 2188 -3196
rect 2132 -3234 2188 -3232
rect 2132 -3286 2134 -3234
rect 2134 -3286 2186 -3234
rect 2186 -3286 2188 -3234
rect 2132 -3288 2188 -3286
rect 2132 -3324 2188 -3322
rect 2132 -3376 2134 -3324
rect 2134 -3376 2186 -3324
rect 2186 -3376 2188 -3324
rect 2132 -3378 2188 -3376
rect 2132 -3414 2188 -3412
rect 2132 -3466 2134 -3414
rect 2134 -3466 2186 -3414
rect 2186 -3466 2188 -3414
rect 2132 -3468 2188 -3466
rect 2132 -3504 2188 -3502
rect 2132 -3556 2134 -3504
rect 2134 -3556 2186 -3504
rect 2186 -3556 2188 -3504
rect 2132 -3558 2188 -3556
rect 2512 -3054 2568 -3052
rect 2512 -3106 2514 -3054
rect 2514 -3106 2566 -3054
rect 2566 -3106 2568 -3054
rect 2512 -3108 2568 -3106
rect 2512 -3144 2568 -3142
rect 2512 -3196 2514 -3144
rect 2514 -3196 2566 -3144
rect 2566 -3196 2568 -3144
rect 2512 -3198 2568 -3196
rect 2512 -3234 2568 -3232
rect 2512 -3286 2514 -3234
rect 2514 -3286 2566 -3234
rect 2566 -3286 2568 -3234
rect 2512 -3288 2568 -3286
rect 2512 -3324 2568 -3322
rect 2512 -3376 2514 -3324
rect 2514 -3376 2566 -3324
rect 2566 -3376 2568 -3324
rect 2512 -3378 2568 -3376
rect 2512 -3414 2568 -3412
rect 2512 -3466 2514 -3414
rect 2514 -3466 2566 -3414
rect 2566 -3466 2568 -3414
rect 2512 -3468 2568 -3466
rect 2512 -3504 2568 -3502
rect 2512 -3556 2514 -3504
rect 2514 -3556 2566 -3504
rect 2566 -3556 2568 -3504
rect 2512 -3558 2568 -3556
rect 2892 -3054 2948 -3052
rect 2892 -3106 2894 -3054
rect 2894 -3106 2946 -3054
rect 2946 -3106 2948 -3054
rect 2892 -3108 2948 -3106
rect 2892 -3144 2948 -3142
rect 2892 -3196 2894 -3144
rect 2894 -3196 2946 -3144
rect 2946 -3196 2948 -3144
rect 2892 -3198 2948 -3196
rect 2892 -3234 2948 -3232
rect 2892 -3286 2894 -3234
rect 2894 -3286 2946 -3234
rect 2946 -3286 2948 -3234
rect 2892 -3288 2948 -3286
rect 2892 -3324 2948 -3322
rect 2892 -3376 2894 -3324
rect 2894 -3376 2946 -3324
rect 2946 -3376 2948 -3324
rect 2892 -3378 2948 -3376
rect 2892 -3414 2948 -3412
rect 2892 -3466 2894 -3414
rect 2894 -3466 2946 -3414
rect 2946 -3466 2948 -3414
rect 2892 -3468 2948 -3466
rect 2892 -3504 2948 -3502
rect 2892 -3556 2894 -3504
rect 2894 -3556 2946 -3504
rect 2946 -3556 2948 -3504
rect 2892 -3558 2948 -3556
rect 3272 -3054 3328 -3052
rect 3272 -3106 3274 -3054
rect 3274 -3106 3326 -3054
rect 3326 -3106 3328 -3054
rect 3272 -3108 3328 -3106
rect 3272 -3144 3328 -3142
rect 3272 -3196 3274 -3144
rect 3274 -3196 3326 -3144
rect 3326 -3196 3328 -3144
rect 3272 -3198 3328 -3196
rect 3272 -3234 3328 -3232
rect 3272 -3286 3274 -3234
rect 3274 -3286 3326 -3234
rect 3326 -3286 3328 -3234
rect 3272 -3288 3328 -3286
rect 3272 -3324 3328 -3322
rect 3272 -3376 3274 -3324
rect 3274 -3376 3326 -3324
rect 3326 -3376 3328 -3324
rect 3272 -3378 3328 -3376
rect 3272 -3414 3328 -3412
rect 3272 -3466 3274 -3414
rect 3274 -3466 3326 -3414
rect 3326 -3466 3328 -3414
rect 3272 -3468 3328 -3466
rect 3272 -3504 3328 -3502
rect 3272 -3556 3274 -3504
rect 3274 -3556 3326 -3504
rect 3326 -3556 3328 -3504
rect 3272 -3558 3328 -3556
rect 3652 -3054 3708 -3052
rect 3652 -3106 3654 -3054
rect 3654 -3106 3706 -3054
rect 3706 -3106 3708 -3054
rect 3652 -3108 3708 -3106
rect 3652 -3144 3708 -3142
rect 3652 -3196 3654 -3144
rect 3654 -3196 3706 -3144
rect 3706 -3196 3708 -3144
rect 3652 -3198 3708 -3196
rect 3652 -3234 3708 -3232
rect 3652 -3286 3654 -3234
rect 3654 -3286 3706 -3234
rect 3706 -3286 3708 -3234
rect 3652 -3288 3708 -3286
rect 3652 -3324 3708 -3322
rect 3652 -3376 3654 -3324
rect 3654 -3376 3706 -3324
rect 3706 -3376 3708 -3324
rect 3652 -3378 3708 -3376
rect 3652 -3414 3708 -3412
rect 3652 -3466 3654 -3414
rect 3654 -3466 3706 -3414
rect 3706 -3466 3708 -3414
rect 3652 -3468 3708 -3466
rect 3652 -3504 3708 -3502
rect 3652 -3556 3654 -3504
rect 3654 -3556 3706 -3504
rect 3706 -3556 3708 -3504
rect 3652 -3558 3708 -3556
rect 4032 -3054 4088 -3052
rect 4032 -3106 4034 -3054
rect 4034 -3106 4086 -3054
rect 4086 -3106 4088 -3054
rect 4032 -3108 4088 -3106
rect 4032 -3144 4088 -3142
rect 4032 -3196 4034 -3144
rect 4034 -3196 4086 -3144
rect 4086 -3196 4088 -3144
rect 4032 -3198 4088 -3196
rect 4032 -3234 4088 -3232
rect 4032 -3286 4034 -3234
rect 4034 -3286 4086 -3234
rect 4086 -3286 4088 -3234
rect 4032 -3288 4088 -3286
rect 4032 -3324 4088 -3322
rect 4032 -3376 4034 -3324
rect 4034 -3376 4086 -3324
rect 4086 -3376 4088 -3324
rect 4032 -3378 4088 -3376
rect 4032 -3414 4088 -3412
rect 4032 -3466 4034 -3414
rect 4034 -3466 4086 -3414
rect 4086 -3466 4088 -3414
rect 4032 -3468 4088 -3466
rect 4032 -3504 4088 -3502
rect 4032 -3556 4034 -3504
rect 4034 -3556 4086 -3504
rect 4086 -3556 4088 -3504
rect 4032 -3558 4088 -3556
rect 4792 -3054 4848 -3052
rect 4792 -3106 4794 -3054
rect 4794 -3106 4846 -3054
rect 4846 -3106 4848 -3054
rect 4792 -3108 4848 -3106
rect 4792 -3144 4848 -3142
rect 4792 -3196 4794 -3144
rect 4794 -3196 4846 -3144
rect 4846 -3196 4848 -3144
rect 4792 -3198 4848 -3196
rect 4792 -3234 4848 -3232
rect 4792 -3286 4794 -3234
rect 4794 -3286 4846 -3234
rect 4846 -3286 4848 -3234
rect 4792 -3288 4848 -3286
rect 4792 -3324 4848 -3322
rect 4792 -3376 4794 -3324
rect 4794 -3376 4846 -3324
rect 4846 -3376 4848 -3324
rect 4792 -3378 4848 -3376
rect 4792 -3414 4848 -3412
rect 4792 -3466 4794 -3414
rect 4794 -3466 4846 -3414
rect 4846 -3466 4848 -3414
rect 4792 -3468 4848 -3466
rect 4792 -3504 4848 -3502
rect 4792 -3556 4794 -3504
rect 4794 -3556 4846 -3504
rect 4846 -3556 4848 -3504
rect 4792 -3558 4848 -3556
rect 5172 -3054 5228 -3052
rect 5172 -3106 5174 -3054
rect 5174 -3106 5226 -3054
rect 5226 -3106 5228 -3054
rect 5172 -3108 5228 -3106
rect 5172 -3144 5228 -3142
rect 5172 -3196 5174 -3144
rect 5174 -3196 5226 -3144
rect 5226 -3196 5228 -3144
rect 5172 -3198 5228 -3196
rect 5172 -3234 5228 -3232
rect 5172 -3286 5174 -3234
rect 5174 -3286 5226 -3234
rect 5226 -3286 5228 -3234
rect 5172 -3288 5228 -3286
rect 5172 -3324 5228 -3322
rect 5172 -3376 5174 -3324
rect 5174 -3376 5226 -3324
rect 5226 -3376 5228 -3324
rect 5172 -3378 5228 -3376
rect 5172 -3414 5228 -3412
rect 5172 -3466 5174 -3414
rect 5174 -3466 5226 -3414
rect 5226 -3466 5228 -3414
rect 5172 -3468 5228 -3466
rect 5172 -3504 5228 -3502
rect 5172 -3556 5174 -3504
rect 5174 -3556 5226 -3504
rect 5226 -3556 5228 -3504
rect 5172 -3558 5228 -3556
rect 5552 -3054 5608 -3052
rect 5552 -3106 5554 -3054
rect 5554 -3106 5606 -3054
rect 5606 -3106 5608 -3054
rect 5552 -3108 5608 -3106
rect 5552 -3144 5608 -3142
rect 5552 -3196 5554 -3144
rect 5554 -3196 5606 -3144
rect 5606 -3196 5608 -3144
rect 5552 -3198 5608 -3196
rect 5552 -3234 5608 -3232
rect 5552 -3286 5554 -3234
rect 5554 -3286 5606 -3234
rect 5606 -3286 5608 -3234
rect 5552 -3288 5608 -3286
rect 5552 -3324 5608 -3322
rect 5552 -3376 5554 -3324
rect 5554 -3376 5606 -3324
rect 5606 -3376 5608 -3324
rect 5552 -3378 5608 -3376
rect 5552 -3414 5608 -3412
rect 5552 -3466 5554 -3414
rect 5554 -3466 5606 -3414
rect 5606 -3466 5608 -3414
rect 5552 -3468 5608 -3466
rect 5552 -3504 5608 -3502
rect 5552 -3556 5554 -3504
rect 5554 -3556 5606 -3504
rect 5606 -3556 5608 -3504
rect 5552 -3558 5608 -3556
rect 5932 -3054 5988 -3052
rect 5932 -3106 5934 -3054
rect 5934 -3106 5986 -3054
rect 5986 -3106 5988 -3054
rect 5932 -3108 5988 -3106
rect 5932 -3144 5988 -3142
rect 5932 -3196 5934 -3144
rect 5934 -3196 5986 -3144
rect 5986 -3196 5988 -3144
rect 5932 -3198 5988 -3196
rect 5932 -3234 5988 -3232
rect 5932 -3286 5934 -3234
rect 5934 -3286 5986 -3234
rect 5986 -3286 5988 -3234
rect 5932 -3288 5988 -3286
rect 5932 -3324 5988 -3322
rect 5932 -3376 5934 -3324
rect 5934 -3376 5986 -3324
rect 5986 -3376 5988 -3324
rect 5932 -3378 5988 -3376
rect 5932 -3414 5988 -3412
rect 5932 -3466 5934 -3414
rect 5934 -3466 5986 -3414
rect 5986 -3466 5988 -3414
rect 5932 -3468 5988 -3466
rect 5932 -3504 5988 -3502
rect 5932 -3556 5934 -3504
rect 5934 -3556 5986 -3504
rect 5986 -3556 5988 -3504
rect 5932 -3558 5988 -3556
rect 6312 -3054 6368 -3052
rect 6312 -3106 6314 -3054
rect 6314 -3106 6366 -3054
rect 6366 -3106 6368 -3054
rect 6312 -3108 6368 -3106
rect 6312 -3144 6368 -3142
rect 6312 -3196 6314 -3144
rect 6314 -3196 6366 -3144
rect 6366 -3196 6368 -3144
rect 6312 -3198 6368 -3196
rect 6312 -3234 6368 -3232
rect 6312 -3286 6314 -3234
rect 6314 -3286 6366 -3234
rect 6366 -3286 6368 -3234
rect 6312 -3288 6368 -3286
rect 6312 -3324 6368 -3322
rect 6312 -3376 6314 -3324
rect 6314 -3376 6366 -3324
rect 6366 -3376 6368 -3324
rect 6312 -3378 6368 -3376
rect 6312 -3414 6368 -3412
rect 6312 -3466 6314 -3414
rect 6314 -3466 6366 -3414
rect 6366 -3466 6368 -3414
rect 6312 -3468 6368 -3466
rect 6312 -3504 6368 -3502
rect 6312 -3556 6314 -3504
rect 6314 -3556 6366 -3504
rect 6366 -3556 6368 -3504
rect 6312 -3558 6368 -3556
rect 6692 -3054 6748 -3052
rect 6692 -3106 6694 -3054
rect 6694 -3106 6746 -3054
rect 6746 -3106 6748 -3054
rect 6692 -3108 6748 -3106
rect 6692 -3144 6748 -3142
rect 6692 -3196 6694 -3144
rect 6694 -3196 6746 -3144
rect 6746 -3196 6748 -3144
rect 6692 -3198 6748 -3196
rect 6692 -3234 6748 -3232
rect 6692 -3286 6694 -3234
rect 6694 -3286 6746 -3234
rect 6746 -3286 6748 -3234
rect 6692 -3288 6748 -3286
rect 6692 -3324 6748 -3322
rect 6692 -3376 6694 -3324
rect 6694 -3376 6746 -3324
rect 6746 -3376 6748 -3324
rect 6692 -3378 6748 -3376
rect 6692 -3414 6748 -3412
rect 6692 -3466 6694 -3414
rect 6694 -3466 6746 -3414
rect 6746 -3466 6748 -3414
rect 6692 -3468 6748 -3466
rect 6692 -3504 6748 -3502
rect 6692 -3556 6694 -3504
rect 6694 -3556 6746 -3504
rect 6746 -3556 6748 -3504
rect 6692 -3558 6748 -3556
rect 7072 -3054 7128 -3052
rect 7072 -3106 7074 -3054
rect 7074 -3106 7126 -3054
rect 7126 -3106 7128 -3054
rect 7072 -3108 7128 -3106
rect 7072 -3144 7128 -3142
rect 7072 -3196 7074 -3144
rect 7074 -3196 7126 -3144
rect 7126 -3196 7128 -3144
rect 7072 -3198 7128 -3196
rect 7072 -3234 7128 -3232
rect 7072 -3286 7074 -3234
rect 7074 -3286 7126 -3234
rect 7126 -3286 7128 -3234
rect 7072 -3288 7128 -3286
rect 7072 -3324 7128 -3322
rect 7072 -3376 7074 -3324
rect 7074 -3376 7126 -3324
rect 7126 -3376 7128 -3324
rect 7072 -3378 7128 -3376
rect 7072 -3414 7128 -3412
rect 7072 -3466 7074 -3414
rect 7074 -3466 7126 -3414
rect 7126 -3466 7128 -3414
rect 7072 -3468 7128 -3466
rect 7072 -3504 7128 -3502
rect 7072 -3556 7074 -3504
rect 7074 -3556 7126 -3504
rect 7126 -3556 7128 -3504
rect 7072 -3558 7128 -3556
rect 7452 -3054 7508 -3052
rect 7452 -3106 7454 -3054
rect 7454 -3106 7506 -3054
rect 7506 -3106 7508 -3054
rect 7452 -3108 7508 -3106
rect 7452 -3144 7508 -3142
rect 7452 -3196 7454 -3144
rect 7454 -3196 7506 -3144
rect 7506 -3196 7508 -3144
rect 7452 -3198 7508 -3196
rect 7452 -3234 7508 -3232
rect 7452 -3286 7454 -3234
rect 7454 -3286 7506 -3234
rect 7506 -3286 7508 -3234
rect 7452 -3288 7508 -3286
rect 7452 -3324 7508 -3322
rect 7452 -3376 7454 -3324
rect 7454 -3376 7506 -3324
rect 7506 -3376 7508 -3324
rect 7452 -3378 7508 -3376
rect 7452 -3414 7508 -3412
rect 7452 -3466 7454 -3414
rect 7454 -3466 7506 -3414
rect 7506 -3466 7508 -3414
rect 7452 -3468 7508 -3466
rect 7452 -3504 7508 -3502
rect 7452 -3556 7454 -3504
rect 7454 -3556 7506 -3504
rect 7506 -3556 7508 -3504
rect 7452 -3558 7508 -3556
rect 7832 -3054 7888 -3052
rect 7832 -3106 7834 -3054
rect 7834 -3106 7886 -3054
rect 7886 -3106 7888 -3054
rect 7832 -3108 7888 -3106
rect 7832 -3144 7888 -3142
rect 7832 -3196 7834 -3144
rect 7834 -3196 7886 -3144
rect 7886 -3196 7888 -3144
rect 7832 -3198 7888 -3196
rect 7832 -3234 7888 -3232
rect 7832 -3286 7834 -3234
rect 7834 -3286 7886 -3234
rect 7886 -3286 7888 -3234
rect 7832 -3288 7888 -3286
rect 7832 -3324 7888 -3322
rect 7832 -3376 7834 -3324
rect 7834 -3376 7886 -3324
rect 7886 -3376 7888 -3324
rect 7832 -3378 7888 -3376
rect 7832 -3414 7888 -3412
rect 7832 -3466 7834 -3414
rect 7834 -3466 7886 -3414
rect 7886 -3466 7888 -3414
rect 7832 -3468 7888 -3466
rect 7832 -3504 7888 -3502
rect 7832 -3556 7834 -3504
rect 7834 -3556 7886 -3504
rect 7886 -3556 7888 -3504
rect 7832 -3558 7888 -3556
rect 8212 -3054 8268 -3052
rect 8212 -3106 8214 -3054
rect 8214 -3106 8266 -3054
rect 8266 -3106 8268 -3054
rect 8212 -3108 8268 -3106
rect 8212 -3144 8268 -3142
rect 8212 -3196 8214 -3144
rect 8214 -3196 8266 -3144
rect 8266 -3196 8268 -3144
rect 8212 -3198 8268 -3196
rect 8212 -3234 8268 -3232
rect 8212 -3286 8214 -3234
rect 8214 -3286 8266 -3234
rect 8266 -3286 8268 -3234
rect 8212 -3288 8268 -3286
rect 8212 -3324 8268 -3322
rect 8212 -3376 8214 -3324
rect 8214 -3376 8266 -3324
rect 8266 -3376 8268 -3324
rect 8212 -3378 8268 -3376
rect 8212 -3414 8268 -3412
rect 8212 -3466 8214 -3414
rect 8214 -3466 8266 -3414
rect 8266 -3466 8268 -3414
rect 8212 -3468 8268 -3466
rect 8212 -3504 8268 -3502
rect 8212 -3556 8214 -3504
rect 8214 -3556 8266 -3504
rect 8266 -3556 8268 -3504
rect 8212 -3558 8268 -3556
rect 4032 -4346 4076 -4302
rect 4076 -4346 4088 -4302
rect 4032 -4358 4088 -4346
rect 4122 -4346 4124 -4302
rect 4124 -4346 4176 -4302
rect 4176 -4346 4178 -4302
rect 4122 -4358 4178 -4346
rect 6312 -4346 6314 -4302
rect 6314 -4346 6366 -4302
rect 6366 -4346 6368 -4302
rect 6312 -4358 6368 -4346
rect 6402 -4346 6404 -4302
rect 6404 -4346 6456 -4302
rect 6456 -4346 6458 -4302
rect 6402 -4358 6458 -4346
rect 8842 -4718 8898 -4662
rect -568 -4828 -512 -4772
rect 8842 -4808 8898 -4752
rect 4032 -4918 4088 -4862
rect 4122 -4918 4178 -4862
rect 4412 -4918 4468 -4862
rect 4502 -4918 4558 -4862
rect -568 -5028 -512 -4972
rect 232 -5028 288 -4972
rect 322 -5028 378 -4972
rect 6312 -5028 6368 -4972
rect 6402 -5028 6458 -4972
rect -98 -5138 -42 -5082
rect -8 -5138 48 -5082
rect -568 -5228 -512 -5172
<< metal3 >>
rect 530 5222 750 5240
rect 530 5158 548 5222
rect 612 5158 668 5222
rect 732 5158 750 5222
rect 530 5140 750 5158
rect 910 5222 1130 5240
rect 910 5158 928 5222
rect 992 5158 1048 5222
rect 1112 5158 1130 5222
rect 910 5140 1130 5158
rect 1290 5222 1510 5240
rect 1290 5158 1308 5222
rect 1372 5158 1428 5222
rect 1492 5158 1510 5222
rect 1290 5140 1510 5158
rect 1670 5222 1890 5240
rect 1670 5158 1688 5222
rect 1752 5158 1808 5222
rect 1872 5158 1890 5222
rect 1670 5140 1890 5158
rect 2050 5222 2270 5240
rect 2050 5158 2068 5222
rect 2132 5158 2188 5222
rect 2252 5158 2270 5222
rect 2050 5140 2270 5158
rect 2430 5222 2650 5240
rect 2430 5158 2448 5222
rect 2512 5158 2568 5222
rect 2632 5158 2650 5222
rect 2430 5140 2650 5158
rect 2810 5222 3030 5240
rect 2810 5158 2828 5222
rect 2892 5158 2948 5222
rect 3012 5158 3030 5222
rect 2810 5140 3030 5158
rect 3190 5222 3410 5240
rect 3190 5158 3208 5222
rect 3272 5158 3328 5222
rect 3392 5158 3410 5222
rect 3190 5140 3410 5158
rect 3570 5222 3790 5240
rect 3570 5158 3588 5222
rect 3652 5158 3708 5222
rect 3772 5158 3790 5222
rect 3570 5140 3790 5158
rect 3950 5222 4170 5240
rect 3950 5158 3968 5222
rect 4032 5158 4088 5222
rect 4152 5158 4170 5222
rect 3950 5140 4170 5158
rect -250 5088 -80 5100
rect -250 5032 -238 5088
rect -182 5032 -148 5088
rect -92 5032 -80 5088
rect -250 5020 -80 5032
rect -250 48 -170 5020
rect -110 4868 60 4880
rect -110 4812 -98 4868
rect -42 4812 -8 4868
rect 48 4812 60 4868
rect -110 4800 60 4812
rect -110 4298 -30 4800
rect -110 4242 -98 4298
rect -42 4242 -30 4298
rect -110 4208 -30 4242
rect -110 4152 -98 4208
rect -42 4152 -30 4208
rect -110 2118 -30 4152
rect -110 2062 -98 2118
rect -42 2062 -30 2118
rect -110 2028 -30 2062
rect -110 1972 -98 2028
rect -42 1972 -30 2028
rect -110 1960 -30 1972
rect 220 4758 390 4770
rect 220 4702 232 4758
rect 288 4702 322 4758
rect 378 4702 390 4758
rect 220 4690 390 4702
rect -250 -8 -238 48
rect -182 -8 -170 48
rect -250 -42 -170 -8
rect -250 -98 -238 -42
rect -182 -98 -170 -42
rect -590 -2112 -490 -2090
rect -590 -2168 -568 -2112
rect -512 -2168 -490 -2112
rect -590 -2190 -490 -2168
rect -250 -2242 -170 -98
rect -250 -2298 -238 -2242
rect -182 -2298 -170 -2242
rect -250 -2332 -170 -2298
rect -250 -2388 -238 -2332
rect -182 -2388 -170 -2332
rect -250 -2400 -170 -2388
rect -110 1798 -30 1820
rect -110 1742 -98 1798
rect -42 1742 -30 1798
rect -110 1708 -30 1742
rect -110 1652 -98 1708
rect -42 1652 -30 1708
rect -110 168 -30 1652
rect -110 112 -98 168
rect -42 112 -30 168
rect -110 78 -30 112
rect -110 22 -98 78
rect -42 22 -30 78
rect -590 -4772 -490 -4750
rect -590 -4828 -568 -4772
rect -512 -4828 -490 -4772
rect -590 -4850 -490 -4828
rect -590 -4972 -490 -4950
rect -590 -5028 -568 -4972
rect -512 -5028 -490 -4972
rect -590 -5050 -490 -5028
rect -110 -5070 -30 22
rect 220 -4960 300 4690
rect 600 3528 680 5140
rect 600 3472 612 3528
rect 668 3472 680 3528
rect 600 3438 680 3472
rect 600 3382 612 3438
rect 668 3382 680 3438
rect 600 3348 680 3382
rect 600 3292 612 3348
rect 668 3292 680 3348
rect 600 3258 680 3292
rect 600 3202 612 3258
rect 668 3202 680 3258
rect 600 3168 680 3202
rect 600 3112 612 3168
rect 668 3112 680 3168
rect 600 3078 680 3112
rect 600 3022 612 3078
rect 668 3022 680 3078
rect 600 1378 680 3022
rect 600 1322 612 1378
rect 668 1322 680 1378
rect 600 1288 680 1322
rect 600 1232 612 1288
rect 668 1232 680 1288
rect 600 1198 680 1232
rect 600 1142 612 1198
rect 668 1142 680 1198
rect 600 1108 680 1142
rect 600 1052 612 1108
rect 668 1052 680 1108
rect 600 1018 680 1052
rect 600 962 612 1018
rect 668 962 680 1018
rect 600 928 680 962
rect 600 872 612 928
rect 668 872 680 928
rect 600 -862 680 872
rect 600 -918 612 -862
rect 668 -918 680 -862
rect 600 -952 680 -918
rect 600 -1008 612 -952
rect 668 -1008 680 -952
rect 600 -1042 680 -1008
rect 600 -1098 612 -1042
rect 668 -1098 680 -1042
rect 600 -1132 680 -1098
rect 600 -1188 612 -1132
rect 668 -1188 680 -1132
rect 600 -1222 680 -1188
rect 600 -1278 612 -1222
rect 668 -1278 680 -1222
rect 600 -1312 680 -1278
rect 600 -1368 612 -1312
rect 668 -1368 680 -1312
rect 600 -3052 680 -1368
rect 600 -3108 612 -3052
rect 668 -3108 680 -3052
rect 600 -3142 680 -3108
rect 600 -3198 612 -3142
rect 668 -3198 680 -3142
rect 600 -3232 680 -3198
rect 600 -3288 612 -3232
rect 668 -3288 680 -3232
rect 600 -3322 680 -3288
rect 600 -3378 612 -3322
rect 668 -3378 680 -3322
rect 600 -3412 680 -3378
rect 600 -3468 612 -3412
rect 668 -3468 680 -3412
rect 600 -3502 680 -3468
rect 600 -3558 612 -3502
rect 668 -3558 680 -3502
rect 600 -4000 680 -3558
rect 980 3528 1060 5140
rect 980 3472 992 3528
rect 1048 3472 1060 3528
rect 980 3438 1060 3472
rect 980 3382 992 3438
rect 1048 3382 1060 3438
rect 980 3348 1060 3382
rect 980 3292 992 3348
rect 1048 3292 1060 3348
rect 980 3258 1060 3292
rect 980 3202 992 3258
rect 1048 3202 1060 3258
rect 980 3168 1060 3202
rect 980 3112 992 3168
rect 1048 3112 1060 3168
rect 980 3078 1060 3112
rect 980 3022 992 3078
rect 1048 3022 1060 3078
rect 980 1378 1060 3022
rect 980 1322 992 1378
rect 1048 1322 1060 1378
rect 980 1288 1060 1322
rect 980 1232 992 1288
rect 1048 1232 1060 1288
rect 980 1198 1060 1232
rect 980 1142 992 1198
rect 1048 1142 1060 1198
rect 980 1108 1060 1142
rect 980 1052 992 1108
rect 1048 1052 1060 1108
rect 980 1018 1060 1052
rect 980 962 992 1018
rect 1048 962 1060 1018
rect 980 928 1060 962
rect 980 872 992 928
rect 1048 872 1060 928
rect 980 -862 1060 872
rect 980 -918 992 -862
rect 1048 -918 1060 -862
rect 980 -952 1060 -918
rect 980 -1008 992 -952
rect 1048 -1008 1060 -952
rect 980 -1042 1060 -1008
rect 980 -1098 992 -1042
rect 1048 -1098 1060 -1042
rect 980 -1132 1060 -1098
rect 980 -1188 992 -1132
rect 1048 -1188 1060 -1132
rect 980 -1222 1060 -1188
rect 980 -1278 992 -1222
rect 1048 -1278 1060 -1222
rect 980 -1312 1060 -1278
rect 980 -1368 992 -1312
rect 1048 -1368 1060 -1312
rect 980 -3052 1060 -1368
rect 980 -3108 992 -3052
rect 1048 -3108 1060 -3052
rect 980 -3142 1060 -3108
rect 980 -3198 992 -3142
rect 1048 -3198 1060 -3142
rect 980 -3232 1060 -3198
rect 980 -3288 992 -3232
rect 1048 -3288 1060 -3232
rect 980 -3322 1060 -3288
rect 980 -3378 992 -3322
rect 1048 -3378 1060 -3322
rect 980 -3412 1060 -3378
rect 980 -3468 992 -3412
rect 1048 -3468 1060 -3412
rect 980 -3502 1060 -3468
rect 980 -3558 992 -3502
rect 1048 -3558 1060 -3502
rect 980 -4000 1060 -3558
rect 1360 3528 1440 5140
rect 1360 3472 1372 3528
rect 1428 3472 1440 3528
rect 1360 3438 1440 3472
rect 1360 3382 1372 3438
rect 1428 3382 1440 3438
rect 1360 3348 1440 3382
rect 1360 3292 1372 3348
rect 1428 3292 1440 3348
rect 1360 3258 1440 3292
rect 1360 3202 1372 3258
rect 1428 3202 1440 3258
rect 1360 3168 1440 3202
rect 1360 3112 1372 3168
rect 1428 3112 1440 3168
rect 1360 3078 1440 3112
rect 1360 3022 1372 3078
rect 1428 3022 1440 3078
rect 1360 1378 1440 3022
rect 1360 1322 1372 1378
rect 1428 1322 1440 1378
rect 1360 1288 1440 1322
rect 1360 1232 1372 1288
rect 1428 1232 1440 1288
rect 1360 1198 1440 1232
rect 1360 1142 1372 1198
rect 1428 1142 1440 1198
rect 1360 1108 1440 1142
rect 1360 1052 1372 1108
rect 1428 1052 1440 1108
rect 1360 1018 1440 1052
rect 1360 962 1372 1018
rect 1428 962 1440 1018
rect 1360 928 1440 962
rect 1360 872 1372 928
rect 1428 872 1440 928
rect 1360 -862 1440 872
rect 1360 -918 1372 -862
rect 1428 -918 1440 -862
rect 1360 -952 1440 -918
rect 1360 -1008 1372 -952
rect 1428 -1008 1440 -952
rect 1360 -1042 1440 -1008
rect 1360 -1098 1372 -1042
rect 1428 -1098 1440 -1042
rect 1360 -1132 1440 -1098
rect 1360 -1188 1372 -1132
rect 1428 -1188 1440 -1132
rect 1360 -1222 1440 -1188
rect 1360 -1278 1372 -1222
rect 1428 -1278 1440 -1222
rect 1360 -1312 1440 -1278
rect 1360 -1368 1372 -1312
rect 1428 -1368 1440 -1312
rect 1360 -3052 1440 -1368
rect 1360 -3108 1372 -3052
rect 1428 -3108 1440 -3052
rect 1360 -3142 1440 -3108
rect 1360 -3198 1372 -3142
rect 1428 -3198 1440 -3142
rect 1360 -3232 1440 -3198
rect 1360 -3288 1372 -3232
rect 1428 -3288 1440 -3232
rect 1360 -3322 1440 -3288
rect 1360 -3378 1372 -3322
rect 1428 -3378 1440 -3322
rect 1360 -3412 1440 -3378
rect 1360 -3468 1372 -3412
rect 1428 -3468 1440 -3412
rect 1360 -3502 1440 -3468
rect 1360 -3558 1372 -3502
rect 1428 -3558 1440 -3502
rect 1360 -4000 1440 -3558
rect 1740 3528 1820 5140
rect 1740 3472 1752 3528
rect 1808 3472 1820 3528
rect 1740 3438 1820 3472
rect 1740 3382 1752 3438
rect 1808 3382 1820 3438
rect 1740 3348 1820 3382
rect 1740 3292 1752 3348
rect 1808 3292 1820 3348
rect 1740 3258 1820 3292
rect 1740 3202 1752 3258
rect 1808 3202 1820 3258
rect 1740 3168 1820 3202
rect 1740 3112 1752 3168
rect 1808 3112 1820 3168
rect 1740 3078 1820 3112
rect 1740 3022 1752 3078
rect 1808 3022 1820 3078
rect 1740 1378 1820 3022
rect 1740 1322 1752 1378
rect 1808 1322 1820 1378
rect 1740 1288 1820 1322
rect 1740 1232 1752 1288
rect 1808 1232 1820 1288
rect 1740 1198 1820 1232
rect 1740 1142 1752 1198
rect 1808 1142 1820 1198
rect 1740 1108 1820 1142
rect 1740 1052 1752 1108
rect 1808 1052 1820 1108
rect 1740 1018 1820 1052
rect 1740 962 1752 1018
rect 1808 962 1820 1018
rect 1740 928 1820 962
rect 1740 872 1752 928
rect 1808 872 1820 928
rect 1740 -862 1820 872
rect 1740 -918 1752 -862
rect 1808 -918 1820 -862
rect 1740 -952 1820 -918
rect 1740 -1008 1752 -952
rect 1808 -1008 1820 -952
rect 1740 -1042 1820 -1008
rect 1740 -1098 1752 -1042
rect 1808 -1098 1820 -1042
rect 1740 -1132 1820 -1098
rect 1740 -1188 1752 -1132
rect 1808 -1188 1820 -1132
rect 1740 -1222 1820 -1188
rect 1740 -1278 1752 -1222
rect 1808 -1278 1820 -1222
rect 1740 -1312 1820 -1278
rect 1740 -1368 1752 -1312
rect 1808 -1368 1820 -1312
rect 1740 -3052 1820 -1368
rect 1740 -3108 1752 -3052
rect 1808 -3108 1820 -3052
rect 1740 -3142 1820 -3108
rect 1740 -3198 1752 -3142
rect 1808 -3198 1820 -3142
rect 1740 -3232 1820 -3198
rect 1740 -3288 1752 -3232
rect 1808 -3288 1820 -3232
rect 1740 -3322 1820 -3288
rect 1740 -3378 1752 -3322
rect 1808 -3378 1820 -3322
rect 1740 -3412 1820 -3378
rect 1740 -3468 1752 -3412
rect 1808 -3468 1820 -3412
rect 1740 -3502 1820 -3468
rect 1740 -3558 1752 -3502
rect 1808 -3558 1820 -3502
rect 1740 -4000 1820 -3558
rect 2120 3528 2200 5140
rect 2120 3472 2132 3528
rect 2188 3472 2200 3528
rect 2120 3438 2200 3472
rect 2120 3382 2132 3438
rect 2188 3382 2200 3438
rect 2120 3348 2200 3382
rect 2120 3292 2132 3348
rect 2188 3292 2200 3348
rect 2120 3258 2200 3292
rect 2120 3202 2132 3258
rect 2188 3202 2200 3258
rect 2120 3168 2200 3202
rect 2120 3112 2132 3168
rect 2188 3112 2200 3168
rect 2120 3078 2200 3112
rect 2120 3022 2132 3078
rect 2188 3022 2200 3078
rect 2120 1378 2200 3022
rect 2120 1322 2132 1378
rect 2188 1322 2200 1378
rect 2120 1288 2200 1322
rect 2120 1232 2132 1288
rect 2188 1232 2200 1288
rect 2120 1198 2200 1232
rect 2120 1142 2132 1198
rect 2188 1142 2200 1198
rect 2120 1108 2200 1142
rect 2120 1052 2132 1108
rect 2188 1052 2200 1108
rect 2120 1018 2200 1052
rect 2120 962 2132 1018
rect 2188 962 2200 1018
rect 2120 928 2200 962
rect 2120 872 2132 928
rect 2188 872 2200 928
rect 2120 -862 2200 872
rect 2120 -918 2132 -862
rect 2188 -918 2200 -862
rect 2120 -952 2200 -918
rect 2120 -1008 2132 -952
rect 2188 -1008 2200 -952
rect 2120 -1042 2200 -1008
rect 2120 -1098 2132 -1042
rect 2188 -1098 2200 -1042
rect 2120 -1132 2200 -1098
rect 2120 -1188 2132 -1132
rect 2188 -1188 2200 -1132
rect 2120 -1222 2200 -1188
rect 2120 -1278 2132 -1222
rect 2188 -1278 2200 -1222
rect 2120 -1312 2200 -1278
rect 2120 -1368 2132 -1312
rect 2188 -1368 2200 -1312
rect 2120 -3052 2200 -1368
rect 2120 -3108 2132 -3052
rect 2188 -3108 2200 -3052
rect 2120 -3142 2200 -3108
rect 2120 -3198 2132 -3142
rect 2188 -3198 2200 -3142
rect 2120 -3232 2200 -3198
rect 2120 -3288 2132 -3232
rect 2188 -3288 2200 -3232
rect 2120 -3322 2200 -3288
rect 2120 -3378 2132 -3322
rect 2188 -3378 2200 -3322
rect 2120 -3412 2200 -3378
rect 2120 -3468 2132 -3412
rect 2188 -3468 2200 -3412
rect 2120 -3502 2200 -3468
rect 2120 -3558 2132 -3502
rect 2188 -3558 2200 -3502
rect 2120 -4000 2200 -3558
rect 2500 3528 2580 5140
rect 2500 3472 2512 3528
rect 2568 3472 2580 3528
rect 2500 3438 2580 3472
rect 2500 3382 2512 3438
rect 2568 3382 2580 3438
rect 2500 3348 2580 3382
rect 2500 3292 2512 3348
rect 2568 3292 2580 3348
rect 2500 3258 2580 3292
rect 2500 3202 2512 3258
rect 2568 3202 2580 3258
rect 2500 3168 2580 3202
rect 2500 3112 2512 3168
rect 2568 3112 2580 3168
rect 2500 3078 2580 3112
rect 2500 3022 2512 3078
rect 2568 3022 2580 3078
rect 2500 1378 2580 3022
rect 2500 1322 2512 1378
rect 2568 1322 2580 1378
rect 2500 1288 2580 1322
rect 2500 1232 2512 1288
rect 2568 1232 2580 1288
rect 2500 1198 2580 1232
rect 2500 1142 2512 1198
rect 2568 1142 2580 1198
rect 2500 1108 2580 1142
rect 2500 1052 2512 1108
rect 2568 1052 2580 1108
rect 2500 1018 2580 1052
rect 2500 962 2512 1018
rect 2568 962 2580 1018
rect 2500 928 2580 962
rect 2500 872 2512 928
rect 2568 872 2580 928
rect 2500 -862 2580 872
rect 2500 -918 2512 -862
rect 2568 -918 2580 -862
rect 2500 -952 2580 -918
rect 2500 -1008 2512 -952
rect 2568 -1008 2580 -952
rect 2500 -1042 2580 -1008
rect 2500 -1098 2512 -1042
rect 2568 -1098 2580 -1042
rect 2500 -1132 2580 -1098
rect 2500 -1188 2512 -1132
rect 2568 -1188 2580 -1132
rect 2500 -1222 2580 -1188
rect 2500 -1278 2512 -1222
rect 2568 -1278 2580 -1222
rect 2500 -1312 2580 -1278
rect 2500 -1368 2512 -1312
rect 2568 -1368 2580 -1312
rect 2500 -3052 2580 -1368
rect 2500 -3108 2512 -3052
rect 2568 -3108 2580 -3052
rect 2500 -3142 2580 -3108
rect 2500 -3198 2512 -3142
rect 2568 -3198 2580 -3142
rect 2500 -3232 2580 -3198
rect 2500 -3288 2512 -3232
rect 2568 -3288 2580 -3232
rect 2500 -3322 2580 -3288
rect 2500 -3378 2512 -3322
rect 2568 -3378 2580 -3322
rect 2500 -3412 2580 -3378
rect 2500 -3468 2512 -3412
rect 2568 -3468 2580 -3412
rect 2500 -3502 2580 -3468
rect 2500 -3558 2512 -3502
rect 2568 -3558 2580 -3502
rect 2500 -4000 2580 -3558
rect 2880 3528 2960 5140
rect 2880 3472 2892 3528
rect 2948 3472 2960 3528
rect 2880 3438 2960 3472
rect 2880 3382 2892 3438
rect 2948 3382 2960 3438
rect 2880 3348 2960 3382
rect 2880 3292 2892 3348
rect 2948 3292 2960 3348
rect 2880 3258 2960 3292
rect 2880 3202 2892 3258
rect 2948 3202 2960 3258
rect 2880 3168 2960 3202
rect 2880 3112 2892 3168
rect 2948 3112 2960 3168
rect 2880 3078 2960 3112
rect 2880 3022 2892 3078
rect 2948 3022 2960 3078
rect 2880 1378 2960 3022
rect 2880 1322 2892 1378
rect 2948 1322 2960 1378
rect 2880 1288 2960 1322
rect 2880 1232 2892 1288
rect 2948 1232 2960 1288
rect 2880 1198 2960 1232
rect 2880 1142 2892 1198
rect 2948 1142 2960 1198
rect 2880 1108 2960 1142
rect 2880 1052 2892 1108
rect 2948 1052 2960 1108
rect 2880 1018 2960 1052
rect 2880 962 2892 1018
rect 2948 962 2960 1018
rect 2880 928 2960 962
rect 2880 872 2892 928
rect 2948 872 2960 928
rect 2880 -862 2960 872
rect 2880 -918 2892 -862
rect 2948 -918 2960 -862
rect 2880 -952 2960 -918
rect 2880 -1008 2892 -952
rect 2948 -1008 2960 -952
rect 2880 -1042 2960 -1008
rect 2880 -1098 2892 -1042
rect 2948 -1098 2960 -1042
rect 2880 -1132 2960 -1098
rect 2880 -1188 2892 -1132
rect 2948 -1188 2960 -1132
rect 2880 -1222 2960 -1188
rect 2880 -1278 2892 -1222
rect 2948 -1278 2960 -1222
rect 2880 -1312 2960 -1278
rect 2880 -1368 2892 -1312
rect 2948 -1368 2960 -1312
rect 2880 -3052 2960 -1368
rect 2880 -3108 2892 -3052
rect 2948 -3108 2960 -3052
rect 2880 -3142 2960 -3108
rect 2880 -3198 2892 -3142
rect 2948 -3198 2960 -3142
rect 2880 -3232 2960 -3198
rect 2880 -3288 2892 -3232
rect 2948 -3288 2960 -3232
rect 2880 -3322 2960 -3288
rect 2880 -3378 2892 -3322
rect 2948 -3378 2960 -3322
rect 2880 -3412 2960 -3378
rect 2880 -3468 2892 -3412
rect 2948 -3468 2960 -3412
rect 2880 -3502 2960 -3468
rect 2880 -3558 2892 -3502
rect 2948 -3558 2960 -3502
rect 2880 -4000 2960 -3558
rect 3260 3528 3340 5140
rect 3260 3472 3272 3528
rect 3328 3472 3340 3528
rect 3260 3438 3340 3472
rect 3260 3382 3272 3438
rect 3328 3382 3340 3438
rect 3260 3348 3340 3382
rect 3260 3292 3272 3348
rect 3328 3292 3340 3348
rect 3260 3258 3340 3292
rect 3260 3202 3272 3258
rect 3328 3202 3340 3258
rect 3260 3168 3340 3202
rect 3260 3112 3272 3168
rect 3328 3112 3340 3168
rect 3260 3078 3340 3112
rect 3260 3022 3272 3078
rect 3328 3022 3340 3078
rect 3260 1378 3340 3022
rect 3260 1322 3272 1378
rect 3328 1322 3340 1378
rect 3260 1288 3340 1322
rect 3260 1232 3272 1288
rect 3328 1232 3340 1288
rect 3260 1198 3340 1232
rect 3260 1142 3272 1198
rect 3328 1142 3340 1198
rect 3260 1108 3340 1142
rect 3260 1052 3272 1108
rect 3328 1052 3340 1108
rect 3260 1018 3340 1052
rect 3260 962 3272 1018
rect 3328 962 3340 1018
rect 3260 928 3340 962
rect 3260 872 3272 928
rect 3328 872 3340 928
rect 3260 -862 3340 872
rect 3260 -918 3272 -862
rect 3328 -918 3340 -862
rect 3260 -952 3340 -918
rect 3260 -1008 3272 -952
rect 3328 -1008 3340 -952
rect 3260 -1042 3340 -1008
rect 3260 -1098 3272 -1042
rect 3328 -1098 3340 -1042
rect 3260 -1132 3340 -1098
rect 3260 -1188 3272 -1132
rect 3328 -1188 3340 -1132
rect 3260 -1222 3340 -1188
rect 3260 -1278 3272 -1222
rect 3328 -1278 3340 -1222
rect 3260 -1312 3340 -1278
rect 3260 -1368 3272 -1312
rect 3328 -1368 3340 -1312
rect 3260 -3052 3340 -1368
rect 3260 -3108 3272 -3052
rect 3328 -3108 3340 -3052
rect 3260 -3142 3340 -3108
rect 3260 -3198 3272 -3142
rect 3328 -3198 3340 -3142
rect 3260 -3232 3340 -3198
rect 3260 -3288 3272 -3232
rect 3328 -3288 3340 -3232
rect 3260 -3322 3340 -3288
rect 3260 -3378 3272 -3322
rect 3328 -3378 3340 -3322
rect 3260 -3412 3340 -3378
rect 3260 -3468 3272 -3412
rect 3328 -3468 3340 -3412
rect 3260 -3502 3340 -3468
rect 3260 -3558 3272 -3502
rect 3328 -3558 3340 -3502
rect 3260 -4000 3340 -3558
rect 3640 3528 3720 5140
rect 3640 3472 3652 3528
rect 3708 3472 3720 3528
rect 3640 3438 3720 3472
rect 3640 3382 3652 3438
rect 3708 3382 3720 3438
rect 3640 3348 3720 3382
rect 3640 3292 3652 3348
rect 3708 3292 3720 3348
rect 3640 3258 3720 3292
rect 3640 3202 3652 3258
rect 3708 3202 3720 3258
rect 3640 3168 3720 3202
rect 3640 3112 3652 3168
rect 3708 3112 3720 3168
rect 3640 3078 3720 3112
rect 3640 3022 3652 3078
rect 3708 3022 3720 3078
rect 3640 1378 3720 3022
rect 3640 1322 3652 1378
rect 3708 1322 3720 1378
rect 3640 1288 3720 1322
rect 3640 1232 3652 1288
rect 3708 1232 3720 1288
rect 3640 1198 3720 1232
rect 3640 1142 3652 1198
rect 3708 1142 3720 1198
rect 3640 1108 3720 1142
rect 3640 1052 3652 1108
rect 3708 1052 3720 1108
rect 3640 1018 3720 1052
rect 3640 962 3652 1018
rect 3708 962 3720 1018
rect 3640 928 3720 962
rect 3640 872 3652 928
rect 3708 872 3720 928
rect 3640 -862 3720 872
rect 3640 -918 3652 -862
rect 3708 -918 3720 -862
rect 3640 -952 3720 -918
rect 3640 -1008 3652 -952
rect 3708 -1008 3720 -952
rect 3640 -1042 3720 -1008
rect 3640 -1098 3652 -1042
rect 3708 -1098 3720 -1042
rect 3640 -1132 3720 -1098
rect 3640 -1188 3652 -1132
rect 3708 -1188 3720 -1132
rect 3640 -1222 3720 -1188
rect 3640 -1278 3652 -1222
rect 3708 -1278 3720 -1222
rect 3640 -1312 3720 -1278
rect 3640 -1368 3652 -1312
rect 3708 -1368 3720 -1312
rect 3640 -3052 3720 -1368
rect 3640 -3108 3652 -3052
rect 3708 -3108 3720 -3052
rect 3640 -3142 3720 -3108
rect 3640 -3198 3652 -3142
rect 3708 -3198 3720 -3142
rect 3640 -3232 3720 -3198
rect 3640 -3288 3652 -3232
rect 3708 -3288 3720 -3232
rect 3640 -3322 3720 -3288
rect 3640 -3378 3652 -3322
rect 3708 -3378 3720 -3322
rect 3640 -3412 3720 -3378
rect 3640 -3468 3652 -3412
rect 3708 -3468 3720 -3412
rect 3640 -3502 3720 -3468
rect 3640 -3558 3652 -3502
rect 3708 -3558 3720 -3502
rect 3640 -4000 3720 -3558
rect 4020 3528 4100 5140
rect 4230 4990 4330 5510
rect 4470 5338 4570 5510
rect 4470 5282 4492 5338
rect 4548 5282 4570 5338
rect 4470 5260 4570 5282
rect 4710 5222 4930 5240
rect 4710 5158 4728 5222
rect 4792 5158 4848 5222
rect 4912 5158 4930 5222
rect 4710 5140 4930 5158
rect 5090 5222 5310 5240
rect 5090 5158 5108 5222
rect 5172 5158 5228 5222
rect 5292 5158 5310 5222
rect 5090 5140 5310 5158
rect 5470 5222 5690 5240
rect 5470 5158 5488 5222
rect 5552 5158 5608 5222
rect 5672 5158 5690 5222
rect 5470 5140 5690 5158
rect 5850 5222 6070 5240
rect 5850 5158 5868 5222
rect 5932 5158 5988 5222
rect 6052 5158 6070 5222
rect 5850 5140 6070 5158
rect 6230 5222 6450 5240
rect 6230 5158 6248 5222
rect 6312 5158 6368 5222
rect 6432 5158 6450 5222
rect 6230 5140 6450 5158
rect 6610 5222 6830 5240
rect 6610 5158 6628 5222
rect 6692 5158 6748 5222
rect 6812 5158 6830 5222
rect 6610 5140 6830 5158
rect 6990 5222 7210 5240
rect 6990 5158 7008 5222
rect 7072 5158 7128 5222
rect 7192 5158 7210 5222
rect 6990 5140 7210 5158
rect 7370 5222 7590 5240
rect 7370 5158 7388 5222
rect 7452 5158 7508 5222
rect 7572 5158 7590 5222
rect 7370 5140 7590 5158
rect 7750 5222 7970 5240
rect 7750 5158 7768 5222
rect 7832 5158 7888 5222
rect 7952 5158 7970 5222
rect 7750 5140 7970 5158
rect 8130 5222 8350 5240
rect 8130 5158 8148 5222
rect 8212 5158 8268 5222
rect 8332 5158 8350 5222
rect 8130 5140 8350 5158
rect 4160 4978 4330 4990
rect 4160 4922 4172 4978
rect 4228 4922 4262 4978
rect 4318 4922 4330 4978
rect 4160 4910 4330 4922
rect 4400 4978 4570 4990
rect 4400 4922 4412 4978
rect 4468 4922 4502 4978
rect 4558 4922 4570 4978
rect 4400 4910 4570 4922
rect 4160 4330 4240 4910
rect 4490 4330 4570 4910
rect 4160 4318 4330 4330
rect 4160 4262 4172 4318
rect 4228 4262 4262 4318
rect 4318 4262 4330 4318
rect 4160 4250 4330 4262
rect 4490 4318 4700 4330
rect 4490 4262 4522 4318
rect 4578 4262 4612 4318
rect 4668 4262 4700 4318
rect 4490 4250 4700 4262
rect 4020 3472 4032 3528
rect 4088 3472 4100 3528
rect 4020 3438 4100 3472
rect 4020 3382 4032 3438
rect 4088 3382 4100 3438
rect 4020 3348 4100 3382
rect 4020 3292 4032 3348
rect 4088 3292 4100 3348
rect 4020 3258 4100 3292
rect 4020 3202 4032 3258
rect 4088 3202 4100 3258
rect 4020 3168 4100 3202
rect 4020 3112 4032 3168
rect 4088 3112 4100 3168
rect 4020 3078 4100 3112
rect 4020 3022 4032 3078
rect 4088 3022 4100 3078
rect 4020 2150 4100 3022
rect 4780 3528 4860 5140
rect 4780 3472 4792 3528
rect 4848 3472 4860 3528
rect 4780 3438 4860 3472
rect 4780 3382 4792 3438
rect 4848 3382 4860 3438
rect 4780 3348 4860 3382
rect 4780 3292 4792 3348
rect 4848 3292 4860 3348
rect 4780 3258 4860 3292
rect 4780 3202 4792 3258
rect 4848 3202 4860 3258
rect 4780 3168 4860 3202
rect 4780 3112 4792 3168
rect 4848 3112 4860 3168
rect 4780 3078 4860 3112
rect 4780 3022 4792 3078
rect 4848 3022 4860 3078
rect 4490 2348 4570 2360
rect 4490 2292 4502 2348
rect 4558 2292 4570 2348
rect 4490 2258 4570 2292
rect 4490 2202 4502 2258
rect 4558 2202 4570 2258
rect 4020 2138 4390 2150
rect 4020 2082 4232 2138
rect 4288 2082 4322 2138
rect 4378 2082 4390 2138
rect 4020 2070 4390 2082
rect 4020 1378 4100 2070
rect 4020 1322 4032 1378
rect 4088 1322 4100 1378
rect 4020 1288 4100 1322
rect 4020 1232 4032 1288
rect 4088 1232 4100 1288
rect 4020 1198 4100 1232
rect 4020 1142 4032 1198
rect 4088 1142 4100 1198
rect 4020 1108 4100 1142
rect 4020 1052 4032 1108
rect 4088 1052 4100 1108
rect 4020 1018 4100 1052
rect 4020 962 4032 1018
rect 4088 962 4100 1018
rect 4020 928 4100 962
rect 4020 872 4032 928
rect 4088 872 4100 928
rect 4020 -862 4100 872
rect 4020 -918 4032 -862
rect 4088 -918 4100 -862
rect 4020 -952 4100 -918
rect 4020 -1008 4032 -952
rect 4088 -1008 4100 -952
rect 4020 -1042 4100 -1008
rect 4020 -1098 4032 -1042
rect 4088 -1098 4100 -1042
rect 4020 -1132 4100 -1098
rect 4020 -1188 4032 -1132
rect 4088 -1188 4100 -1132
rect 4020 -1222 4100 -1188
rect 4020 -1278 4032 -1222
rect 4088 -1278 4100 -1222
rect 4020 -1312 4100 -1278
rect 4020 -1368 4032 -1312
rect 4088 -1368 4100 -1312
rect 4020 -3052 4100 -1368
rect 4020 -3108 4032 -3052
rect 4088 -3108 4100 -3052
rect 4020 -3142 4100 -3108
rect 4020 -3198 4032 -3142
rect 4088 -3198 4100 -3142
rect 4020 -3232 4100 -3198
rect 4020 -3288 4032 -3232
rect 4088 -3288 4100 -3232
rect 4020 -3322 4100 -3288
rect 4020 -3378 4032 -3322
rect 4088 -3378 4100 -3322
rect 4020 -3412 4100 -3378
rect 4020 -3468 4032 -3412
rect 4088 -3468 4100 -3412
rect 4020 -3502 4100 -3468
rect 4020 -3558 4032 -3502
rect 4088 -3558 4100 -3502
rect 4020 -4000 4100 -3558
rect 4490 168 4570 2202
rect 4490 112 4502 168
rect 4558 112 4570 168
rect 4490 78 4570 112
rect 4490 22 4502 78
rect 4558 22 4570 78
rect 4020 -4302 4190 -4290
rect 4020 -4358 4032 -4302
rect 4088 -4358 4122 -4302
rect 4178 -4358 4190 -4302
rect 4020 -4370 4190 -4358
rect 4110 -4850 4190 -4370
rect 4490 -4850 4570 22
rect 4780 1378 4860 3022
rect 4780 1322 4792 1378
rect 4848 1322 4860 1378
rect 4780 1288 4860 1322
rect 4780 1232 4792 1288
rect 4848 1232 4860 1288
rect 4780 1198 4860 1232
rect 4780 1142 4792 1198
rect 4848 1142 4860 1198
rect 4780 1108 4860 1142
rect 4780 1052 4792 1108
rect 4848 1052 4860 1108
rect 4780 1018 4860 1052
rect 4780 962 4792 1018
rect 4848 962 4860 1018
rect 4780 928 4860 962
rect 4780 872 4792 928
rect 4848 872 4860 928
rect 4780 -862 4860 872
rect 4780 -918 4792 -862
rect 4848 -918 4860 -862
rect 4780 -952 4860 -918
rect 4780 -1008 4792 -952
rect 4848 -1008 4860 -952
rect 4780 -1042 4860 -1008
rect 4780 -1098 4792 -1042
rect 4848 -1098 4860 -1042
rect 4780 -1132 4860 -1098
rect 4780 -1188 4792 -1132
rect 4848 -1188 4860 -1132
rect 4780 -1222 4860 -1188
rect 4780 -1278 4792 -1222
rect 4848 -1278 4860 -1222
rect 4780 -1312 4860 -1278
rect 4780 -1368 4792 -1312
rect 4848 -1368 4860 -1312
rect 4780 -3052 4860 -1368
rect 4780 -3108 4792 -3052
rect 4848 -3108 4860 -3052
rect 4780 -3142 4860 -3108
rect 4780 -3198 4792 -3142
rect 4848 -3198 4860 -3142
rect 4780 -3232 4860 -3198
rect 4780 -3288 4792 -3232
rect 4848 -3288 4860 -3232
rect 4780 -3322 4860 -3288
rect 4780 -3378 4792 -3322
rect 4848 -3378 4860 -3322
rect 4780 -3412 4860 -3378
rect 4780 -3468 4792 -3412
rect 4848 -3468 4860 -3412
rect 4780 -3502 4860 -3468
rect 4780 -3558 4792 -3502
rect 4848 -3558 4860 -3502
rect 4780 -4000 4860 -3558
rect 5160 3528 5240 5140
rect 5160 3472 5172 3528
rect 5228 3472 5240 3528
rect 5160 3438 5240 3472
rect 5160 3382 5172 3438
rect 5228 3382 5240 3438
rect 5160 3348 5240 3382
rect 5160 3292 5172 3348
rect 5228 3292 5240 3348
rect 5160 3258 5240 3292
rect 5160 3202 5172 3258
rect 5228 3202 5240 3258
rect 5160 3168 5240 3202
rect 5160 3112 5172 3168
rect 5228 3112 5240 3168
rect 5160 3078 5240 3112
rect 5160 3022 5172 3078
rect 5228 3022 5240 3078
rect 5160 1378 5240 3022
rect 5160 1322 5172 1378
rect 5228 1322 5240 1378
rect 5160 1288 5240 1322
rect 5160 1232 5172 1288
rect 5228 1232 5240 1288
rect 5160 1198 5240 1232
rect 5160 1142 5172 1198
rect 5228 1142 5240 1198
rect 5160 1108 5240 1142
rect 5160 1052 5172 1108
rect 5228 1052 5240 1108
rect 5160 1018 5240 1052
rect 5160 962 5172 1018
rect 5228 962 5240 1018
rect 5160 928 5240 962
rect 5160 872 5172 928
rect 5228 872 5240 928
rect 5160 -862 5240 872
rect 5160 -918 5172 -862
rect 5228 -918 5240 -862
rect 5160 -952 5240 -918
rect 5160 -1008 5172 -952
rect 5228 -1008 5240 -952
rect 5160 -1042 5240 -1008
rect 5160 -1098 5172 -1042
rect 5228 -1098 5240 -1042
rect 5160 -1132 5240 -1098
rect 5160 -1188 5172 -1132
rect 5228 -1188 5240 -1132
rect 5160 -1222 5240 -1188
rect 5160 -1278 5172 -1222
rect 5228 -1278 5240 -1222
rect 5160 -1312 5240 -1278
rect 5160 -1368 5172 -1312
rect 5228 -1368 5240 -1312
rect 5160 -3052 5240 -1368
rect 5160 -3108 5172 -3052
rect 5228 -3108 5240 -3052
rect 5160 -3142 5240 -3108
rect 5160 -3198 5172 -3142
rect 5228 -3198 5240 -3142
rect 5160 -3232 5240 -3198
rect 5160 -3288 5172 -3232
rect 5228 -3288 5240 -3232
rect 5160 -3322 5240 -3288
rect 5160 -3378 5172 -3322
rect 5228 -3378 5240 -3322
rect 5160 -3412 5240 -3378
rect 5160 -3468 5172 -3412
rect 5228 -3468 5240 -3412
rect 5160 -3502 5240 -3468
rect 5160 -3558 5172 -3502
rect 5228 -3558 5240 -3502
rect 5160 -4000 5240 -3558
rect 5540 3528 5620 5140
rect 5540 3472 5552 3528
rect 5608 3472 5620 3528
rect 5540 3438 5620 3472
rect 5540 3382 5552 3438
rect 5608 3382 5620 3438
rect 5540 3348 5620 3382
rect 5540 3292 5552 3348
rect 5608 3292 5620 3348
rect 5540 3258 5620 3292
rect 5540 3202 5552 3258
rect 5608 3202 5620 3258
rect 5540 3168 5620 3202
rect 5540 3112 5552 3168
rect 5608 3112 5620 3168
rect 5540 3078 5620 3112
rect 5540 3022 5552 3078
rect 5608 3022 5620 3078
rect 5540 1378 5620 3022
rect 5540 1322 5552 1378
rect 5608 1322 5620 1378
rect 5540 1288 5620 1322
rect 5540 1232 5552 1288
rect 5608 1232 5620 1288
rect 5540 1198 5620 1232
rect 5540 1142 5552 1198
rect 5608 1142 5620 1198
rect 5540 1108 5620 1142
rect 5540 1052 5552 1108
rect 5608 1052 5620 1108
rect 5540 1018 5620 1052
rect 5540 962 5552 1018
rect 5608 962 5620 1018
rect 5540 928 5620 962
rect 5540 872 5552 928
rect 5608 872 5620 928
rect 5540 -862 5620 872
rect 5540 -918 5552 -862
rect 5608 -918 5620 -862
rect 5540 -952 5620 -918
rect 5540 -1008 5552 -952
rect 5608 -1008 5620 -952
rect 5540 -1042 5620 -1008
rect 5540 -1098 5552 -1042
rect 5608 -1098 5620 -1042
rect 5540 -1132 5620 -1098
rect 5540 -1188 5552 -1132
rect 5608 -1188 5620 -1132
rect 5540 -1222 5620 -1188
rect 5540 -1278 5552 -1222
rect 5608 -1278 5620 -1222
rect 5540 -1312 5620 -1278
rect 5540 -1368 5552 -1312
rect 5608 -1368 5620 -1312
rect 5540 -3052 5620 -1368
rect 5540 -3108 5552 -3052
rect 5608 -3108 5620 -3052
rect 5540 -3142 5620 -3108
rect 5540 -3198 5552 -3142
rect 5608 -3198 5620 -3142
rect 5540 -3232 5620 -3198
rect 5540 -3288 5552 -3232
rect 5608 -3288 5620 -3232
rect 5540 -3322 5620 -3288
rect 5540 -3378 5552 -3322
rect 5608 -3378 5620 -3322
rect 5540 -3412 5620 -3378
rect 5540 -3468 5552 -3412
rect 5608 -3468 5620 -3412
rect 5540 -3502 5620 -3468
rect 5540 -3558 5552 -3502
rect 5608 -3558 5620 -3502
rect 5540 -4000 5620 -3558
rect 5920 3528 6000 5140
rect 5920 3472 5932 3528
rect 5988 3472 6000 3528
rect 5920 3438 6000 3472
rect 5920 3382 5932 3438
rect 5988 3382 6000 3438
rect 5920 3348 6000 3382
rect 5920 3292 5932 3348
rect 5988 3292 6000 3348
rect 5920 3258 6000 3292
rect 5920 3202 5932 3258
rect 5988 3202 6000 3258
rect 5920 3168 6000 3202
rect 5920 3112 5932 3168
rect 5988 3112 6000 3168
rect 5920 3078 6000 3112
rect 5920 3022 5932 3078
rect 5988 3022 6000 3078
rect 5920 1378 6000 3022
rect 5920 1322 5932 1378
rect 5988 1322 6000 1378
rect 5920 1288 6000 1322
rect 5920 1232 5932 1288
rect 5988 1232 6000 1288
rect 5920 1198 6000 1232
rect 5920 1142 5932 1198
rect 5988 1142 6000 1198
rect 5920 1108 6000 1142
rect 5920 1052 5932 1108
rect 5988 1052 6000 1108
rect 5920 1018 6000 1052
rect 5920 962 5932 1018
rect 5988 962 6000 1018
rect 5920 928 6000 962
rect 5920 872 5932 928
rect 5988 872 6000 928
rect 5920 -862 6000 872
rect 5920 -918 5932 -862
rect 5988 -918 6000 -862
rect 5920 -952 6000 -918
rect 5920 -1008 5932 -952
rect 5988 -1008 6000 -952
rect 5920 -1042 6000 -1008
rect 5920 -1098 5932 -1042
rect 5988 -1098 6000 -1042
rect 5920 -1132 6000 -1098
rect 5920 -1188 5932 -1132
rect 5988 -1188 6000 -1132
rect 5920 -1222 6000 -1188
rect 5920 -1278 5932 -1222
rect 5988 -1278 6000 -1222
rect 5920 -1312 6000 -1278
rect 5920 -1368 5932 -1312
rect 5988 -1368 6000 -1312
rect 5920 -3052 6000 -1368
rect 5920 -3108 5932 -3052
rect 5988 -3108 6000 -3052
rect 5920 -3142 6000 -3108
rect 5920 -3198 5932 -3142
rect 5988 -3198 6000 -3142
rect 5920 -3232 6000 -3198
rect 5920 -3288 5932 -3232
rect 5988 -3288 6000 -3232
rect 5920 -3322 6000 -3288
rect 5920 -3378 5932 -3322
rect 5988 -3378 6000 -3322
rect 5920 -3412 6000 -3378
rect 5920 -3468 5932 -3412
rect 5988 -3468 6000 -3412
rect 5920 -3502 6000 -3468
rect 5920 -3558 5932 -3502
rect 5988 -3558 6000 -3502
rect 5920 -4000 6000 -3558
rect 6300 3528 6380 5140
rect 6300 3472 6312 3528
rect 6368 3472 6380 3528
rect 6300 3438 6380 3472
rect 6300 3382 6312 3438
rect 6368 3382 6380 3438
rect 6300 3348 6380 3382
rect 6300 3292 6312 3348
rect 6368 3292 6380 3348
rect 6300 3258 6380 3292
rect 6300 3202 6312 3258
rect 6368 3202 6380 3258
rect 6300 3168 6380 3202
rect 6300 3112 6312 3168
rect 6368 3112 6380 3168
rect 6300 3078 6380 3112
rect 6300 3022 6312 3078
rect 6368 3022 6380 3078
rect 6300 1378 6380 3022
rect 6300 1322 6312 1378
rect 6368 1322 6380 1378
rect 6300 1288 6380 1322
rect 6300 1232 6312 1288
rect 6368 1232 6380 1288
rect 6300 1198 6380 1232
rect 6300 1142 6312 1198
rect 6368 1142 6380 1198
rect 6300 1108 6380 1142
rect 6300 1052 6312 1108
rect 6368 1052 6380 1108
rect 6300 1018 6380 1052
rect 6300 962 6312 1018
rect 6368 962 6380 1018
rect 6300 928 6380 962
rect 6300 872 6312 928
rect 6368 872 6380 928
rect 6300 -862 6380 872
rect 6300 -918 6312 -862
rect 6368 -918 6380 -862
rect 6300 -952 6380 -918
rect 6300 -1008 6312 -952
rect 6368 -1008 6380 -952
rect 6300 -1042 6380 -1008
rect 6300 -1098 6312 -1042
rect 6368 -1098 6380 -1042
rect 6300 -1132 6380 -1098
rect 6300 -1188 6312 -1132
rect 6368 -1188 6380 -1132
rect 6300 -1222 6380 -1188
rect 6300 -1278 6312 -1222
rect 6368 -1278 6380 -1222
rect 6300 -1312 6380 -1278
rect 6300 -1368 6312 -1312
rect 6368 -1368 6380 -1312
rect 6300 -3052 6380 -1368
rect 6300 -3108 6312 -3052
rect 6368 -3108 6380 -3052
rect 6300 -3142 6380 -3108
rect 6300 -3198 6312 -3142
rect 6368 -3198 6380 -3142
rect 6300 -3232 6380 -3198
rect 6300 -3288 6312 -3232
rect 6368 -3288 6380 -3232
rect 6300 -3322 6380 -3288
rect 6300 -3378 6312 -3322
rect 6368 -3378 6380 -3322
rect 6300 -3412 6380 -3378
rect 6300 -3468 6312 -3412
rect 6368 -3468 6380 -3412
rect 6300 -3502 6380 -3468
rect 6300 -3558 6312 -3502
rect 6368 -3558 6380 -3502
rect 6300 -4000 6380 -3558
rect 6680 3528 6760 5140
rect 6680 3472 6692 3528
rect 6748 3472 6760 3528
rect 6680 3438 6760 3472
rect 6680 3382 6692 3438
rect 6748 3382 6760 3438
rect 6680 3348 6760 3382
rect 6680 3292 6692 3348
rect 6748 3292 6760 3348
rect 6680 3258 6760 3292
rect 6680 3202 6692 3258
rect 6748 3202 6760 3258
rect 6680 3168 6760 3202
rect 6680 3112 6692 3168
rect 6748 3112 6760 3168
rect 6680 3078 6760 3112
rect 6680 3022 6692 3078
rect 6748 3022 6760 3078
rect 6680 1378 6760 3022
rect 6680 1322 6692 1378
rect 6748 1322 6760 1378
rect 6680 1288 6760 1322
rect 6680 1232 6692 1288
rect 6748 1232 6760 1288
rect 6680 1198 6760 1232
rect 6680 1142 6692 1198
rect 6748 1142 6760 1198
rect 6680 1108 6760 1142
rect 6680 1052 6692 1108
rect 6748 1052 6760 1108
rect 6680 1018 6760 1052
rect 6680 962 6692 1018
rect 6748 962 6760 1018
rect 6680 928 6760 962
rect 6680 872 6692 928
rect 6748 872 6760 928
rect 6680 -862 6760 872
rect 6680 -918 6692 -862
rect 6748 -918 6760 -862
rect 6680 -952 6760 -918
rect 6680 -1008 6692 -952
rect 6748 -1008 6760 -952
rect 6680 -1042 6760 -1008
rect 6680 -1098 6692 -1042
rect 6748 -1098 6760 -1042
rect 6680 -1132 6760 -1098
rect 6680 -1188 6692 -1132
rect 6748 -1188 6760 -1132
rect 6680 -1222 6760 -1188
rect 6680 -1278 6692 -1222
rect 6748 -1278 6760 -1222
rect 6680 -1312 6760 -1278
rect 6680 -1368 6692 -1312
rect 6748 -1368 6760 -1312
rect 6680 -3052 6760 -1368
rect 6680 -3108 6692 -3052
rect 6748 -3108 6760 -3052
rect 6680 -3142 6760 -3108
rect 6680 -3198 6692 -3142
rect 6748 -3198 6760 -3142
rect 6680 -3232 6760 -3198
rect 6680 -3288 6692 -3232
rect 6748 -3288 6760 -3232
rect 6680 -3322 6760 -3288
rect 6680 -3378 6692 -3322
rect 6748 -3378 6760 -3322
rect 6680 -3412 6760 -3378
rect 6680 -3468 6692 -3412
rect 6748 -3468 6760 -3412
rect 6680 -3502 6760 -3468
rect 6680 -3558 6692 -3502
rect 6748 -3558 6760 -3502
rect 6680 -4000 6760 -3558
rect 7060 3528 7140 5140
rect 7060 3472 7072 3528
rect 7128 3472 7140 3528
rect 7060 3438 7140 3472
rect 7060 3382 7072 3438
rect 7128 3382 7140 3438
rect 7060 3348 7140 3382
rect 7060 3292 7072 3348
rect 7128 3292 7140 3348
rect 7060 3258 7140 3292
rect 7060 3202 7072 3258
rect 7128 3202 7140 3258
rect 7060 3168 7140 3202
rect 7060 3112 7072 3168
rect 7128 3112 7140 3168
rect 7060 3078 7140 3112
rect 7060 3022 7072 3078
rect 7128 3022 7140 3078
rect 7060 1378 7140 3022
rect 7060 1322 7072 1378
rect 7128 1322 7140 1378
rect 7060 1288 7140 1322
rect 7060 1232 7072 1288
rect 7128 1232 7140 1288
rect 7060 1198 7140 1232
rect 7060 1142 7072 1198
rect 7128 1142 7140 1198
rect 7060 1108 7140 1142
rect 7060 1052 7072 1108
rect 7128 1052 7140 1108
rect 7060 1018 7140 1052
rect 7060 962 7072 1018
rect 7128 962 7140 1018
rect 7060 928 7140 962
rect 7060 872 7072 928
rect 7128 872 7140 928
rect 7060 -862 7140 872
rect 7060 -918 7072 -862
rect 7128 -918 7140 -862
rect 7060 -952 7140 -918
rect 7060 -1008 7072 -952
rect 7128 -1008 7140 -952
rect 7060 -1042 7140 -1008
rect 7060 -1098 7072 -1042
rect 7128 -1098 7140 -1042
rect 7060 -1132 7140 -1098
rect 7060 -1188 7072 -1132
rect 7128 -1188 7140 -1132
rect 7060 -1222 7140 -1188
rect 7060 -1278 7072 -1222
rect 7128 -1278 7140 -1222
rect 7060 -1312 7140 -1278
rect 7060 -1368 7072 -1312
rect 7128 -1368 7140 -1312
rect 7060 -3052 7140 -1368
rect 7060 -3108 7072 -3052
rect 7128 -3108 7140 -3052
rect 7060 -3142 7140 -3108
rect 7060 -3198 7072 -3142
rect 7128 -3198 7140 -3142
rect 7060 -3232 7140 -3198
rect 7060 -3288 7072 -3232
rect 7128 -3288 7140 -3232
rect 7060 -3322 7140 -3288
rect 7060 -3378 7072 -3322
rect 7128 -3378 7140 -3322
rect 7060 -3412 7140 -3378
rect 7060 -3468 7072 -3412
rect 7128 -3468 7140 -3412
rect 7060 -3502 7140 -3468
rect 7060 -3558 7072 -3502
rect 7128 -3558 7140 -3502
rect 7060 -4000 7140 -3558
rect 7440 3528 7520 5140
rect 7440 3472 7452 3528
rect 7508 3472 7520 3528
rect 7440 3438 7520 3472
rect 7440 3382 7452 3438
rect 7508 3382 7520 3438
rect 7440 3348 7520 3382
rect 7440 3292 7452 3348
rect 7508 3292 7520 3348
rect 7440 3258 7520 3292
rect 7440 3202 7452 3258
rect 7508 3202 7520 3258
rect 7440 3168 7520 3202
rect 7440 3112 7452 3168
rect 7508 3112 7520 3168
rect 7440 3078 7520 3112
rect 7440 3022 7452 3078
rect 7508 3022 7520 3078
rect 7440 1378 7520 3022
rect 7440 1322 7452 1378
rect 7508 1322 7520 1378
rect 7440 1288 7520 1322
rect 7440 1232 7452 1288
rect 7508 1232 7520 1288
rect 7440 1198 7520 1232
rect 7440 1142 7452 1198
rect 7508 1142 7520 1198
rect 7440 1108 7520 1142
rect 7440 1052 7452 1108
rect 7508 1052 7520 1108
rect 7440 1018 7520 1052
rect 7440 962 7452 1018
rect 7508 962 7520 1018
rect 7440 928 7520 962
rect 7440 872 7452 928
rect 7508 872 7520 928
rect 7440 -862 7520 872
rect 7440 -918 7452 -862
rect 7508 -918 7520 -862
rect 7440 -952 7520 -918
rect 7440 -1008 7452 -952
rect 7508 -1008 7520 -952
rect 7440 -1042 7520 -1008
rect 7440 -1098 7452 -1042
rect 7508 -1098 7520 -1042
rect 7440 -1132 7520 -1098
rect 7440 -1188 7452 -1132
rect 7508 -1188 7520 -1132
rect 7440 -1222 7520 -1188
rect 7440 -1278 7452 -1222
rect 7508 -1278 7520 -1222
rect 7440 -1312 7520 -1278
rect 7440 -1368 7452 -1312
rect 7508 -1368 7520 -1312
rect 7440 -3052 7520 -1368
rect 7440 -3108 7452 -3052
rect 7508 -3108 7520 -3052
rect 7440 -3142 7520 -3108
rect 7440 -3198 7452 -3142
rect 7508 -3198 7520 -3142
rect 7440 -3232 7520 -3198
rect 7440 -3288 7452 -3232
rect 7508 -3288 7520 -3232
rect 7440 -3322 7520 -3288
rect 7440 -3378 7452 -3322
rect 7508 -3378 7520 -3322
rect 7440 -3412 7520 -3378
rect 7440 -3468 7452 -3412
rect 7508 -3468 7520 -3412
rect 7440 -3502 7520 -3468
rect 7440 -3558 7452 -3502
rect 7508 -3558 7520 -3502
rect 7440 -4000 7520 -3558
rect 7820 3528 7900 5140
rect 7820 3472 7832 3528
rect 7888 3472 7900 3528
rect 7820 3438 7900 3472
rect 7820 3382 7832 3438
rect 7888 3382 7900 3438
rect 7820 3348 7900 3382
rect 7820 3292 7832 3348
rect 7888 3292 7900 3348
rect 7820 3258 7900 3292
rect 7820 3202 7832 3258
rect 7888 3202 7900 3258
rect 7820 3168 7900 3202
rect 7820 3112 7832 3168
rect 7888 3112 7900 3168
rect 7820 3078 7900 3112
rect 7820 3022 7832 3078
rect 7888 3022 7900 3078
rect 7820 1378 7900 3022
rect 7820 1322 7832 1378
rect 7888 1322 7900 1378
rect 7820 1288 7900 1322
rect 7820 1232 7832 1288
rect 7888 1232 7900 1288
rect 7820 1198 7900 1232
rect 7820 1142 7832 1198
rect 7888 1142 7900 1198
rect 7820 1108 7900 1142
rect 7820 1052 7832 1108
rect 7888 1052 7900 1108
rect 7820 1018 7900 1052
rect 7820 962 7832 1018
rect 7888 962 7900 1018
rect 7820 928 7900 962
rect 7820 872 7832 928
rect 7888 872 7900 928
rect 7820 -862 7900 872
rect 7820 -918 7832 -862
rect 7888 -918 7900 -862
rect 7820 -952 7900 -918
rect 7820 -1008 7832 -952
rect 7888 -1008 7900 -952
rect 7820 -1042 7900 -1008
rect 7820 -1098 7832 -1042
rect 7888 -1098 7900 -1042
rect 7820 -1132 7900 -1098
rect 7820 -1188 7832 -1132
rect 7888 -1188 7900 -1132
rect 7820 -1222 7900 -1188
rect 7820 -1278 7832 -1222
rect 7888 -1278 7900 -1222
rect 7820 -1312 7900 -1278
rect 7820 -1368 7832 -1312
rect 7888 -1368 7900 -1312
rect 7820 -3052 7900 -1368
rect 7820 -3108 7832 -3052
rect 7888 -3108 7900 -3052
rect 7820 -3142 7900 -3108
rect 7820 -3198 7832 -3142
rect 7888 -3198 7900 -3142
rect 7820 -3232 7900 -3198
rect 7820 -3288 7832 -3232
rect 7888 -3288 7900 -3232
rect 7820 -3322 7900 -3288
rect 7820 -3378 7832 -3322
rect 7888 -3378 7900 -3322
rect 7820 -3412 7900 -3378
rect 7820 -3468 7832 -3412
rect 7888 -3468 7900 -3412
rect 7820 -3502 7900 -3468
rect 7820 -3558 7832 -3502
rect 7888 -3558 7900 -3502
rect 7820 -4000 7900 -3558
rect 8200 3528 8280 5140
rect 8600 4868 8770 4880
rect 8600 4812 8612 4868
rect 8668 4812 8702 4868
rect 8758 4812 8770 4868
rect 8600 4800 8770 4812
rect 8200 3472 8212 3528
rect 8268 3472 8280 3528
rect 8200 3438 8280 3472
rect 8200 3382 8212 3438
rect 8268 3382 8280 3438
rect 8200 3348 8280 3382
rect 8200 3292 8212 3348
rect 8268 3292 8280 3348
rect 8200 3258 8280 3292
rect 8200 3202 8212 3258
rect 8268 3202 8280 3258
rect 8200 3168 8280 3202
rect 8200 3112 8212 3168
rect 8268 3112 8280 3168
rect 8200 3078 8280 3112
rect 8200 3022 8212 3078
rect 8268 3022 8280 3078
rect 8200 1378 8280 3022
rect 8200 1322 8212 1378
rect 8268 1322 8280 1378
rect 8200 1288 8280 1322
rect 8200 1232 8212 1288
rect 8268 1232 8280 1288
rect 8200 1198 8280 1232
rect 8200 1142 8212 1198
rect 8268 1142 8280 1198
rect 8200 1108 8280 1142
rect 8200 1052 8212 1108
rect 8268 1052 8280 1108
rect 8200 1018 8280 1052
rect 8200 962 8212 1018
rect 8268 962 8280 1018
rect 8200 928 8280 962
rect 8200 872 8212 928
rect 8268 872 8280 928
rect 8200 -862 8280 872
rect 8200 -918 8212 -862
rect 8268 -918 8280 -862
rect 8200 -952 8280 -918
rect 8200 -1008 8212 -952
rect 8268 -1008 8280 -952
rect 8200 -1042 8280 -1008
rect 8200 -1098 8212 -1042
rect 8268 -1098 8280 -1042
rect 8200 -1132 8280 -1098
rect 8200 -1188 8212 -1132
rect 8268 -1188 8280 -1132
rect 8200 -1222 8280 -1188
rect 8200 -1278 8212 -1222
rect 8268 -1278 8280 -1222
rect 8200 -1312 8280 -1278
rect 8200 -1368 8212 -1312
rect 8268 -1368 8280 -1312
rect 8200 -3052 8280 -1368
rect 8690 -62 8770 4800
rect 8690 -118 8702 -62
rect 8758 -118 8770 -62
rect 8690 -152 8770 -118
rect 8690 -208 8702 -152
rect 8758 -208 8770 -152
rect 8690 -2242 8770 -208
rect 8690 -2298 8702 -2242
rect 8758 -2298 8770 -2242
rect 8690 -2332 8770 -2298
rect 8690 -2388 8702 -2332
rect 8758 -2388 8770 -2332
rect 8690 -2400 8770 -2388
rect 8830 2348 8910 2370
rect 8830 2292 8842 2348
rect 8898 2292 8910 2348
rect 8830 2258 8910 2292
rect 8830 2202 8842 2258
rect 8898 2202 8910 2258
rect 8830 168 8910 2202
rect 8830 112 8842 168
rect 8898 112 8910 168
rect 8830 78 8910 112
rect 8830 22 8842 78
rect 8898 22 8910 78
rect 8200 -3108 8212 -3052
rect 8268 -3108 8280 -3052
rect 8200 -3142 8280 -3108
rect 8200 -3198 8212 -3142
rect 8268 -3198 8280 -3142
rect 8200 -3232 8280 -3198
rect 8200 -3288 8212 -3232
rect 8268 -3288 8280 -3232
rect 8200 -3322 8280 -3288
rect 8200 -3378 8212 -3322
rect 8268 -3378 8280 -3322
rect 8200 -3412 8280 -3378
rect 8200 -3468 8212 -3412
rect 8268 -3468 8280 -3412
rect 8200 -3502 8280 -3468
rect 8200 -3558 8212 -3502
rect 8268 -3558 8280 -3502
rect 8200 -4000 8280 -3558
rect 6300 -4302 6470 -4290
rect 6300 -4358 6312 -4302
rect 6368 -4358 6402 -4302
rect 6458 -4358 6470 -4302
rect 6300 -4370 6470 -4358
rect 4020 -4862 4190 -4850
rect 4020 -4918 4032 -4862
rect 4088 -4918 4122 -4862
rect 4178 -4918 4190 -4862
rect 4020 -4930 4190 -4918
rect 4400 -4862 4570 -4850
rect 4400 -4918 4412 -4862
rect 4468 -4918 4502 -4862
rect 4558 -4918 4570 -4862
rect 4400 -4930 4570 -4918
rect 6390 -4960 6470 -4370
rect 8830 -4662 8910 22
rect 8830 -4718 8842 -4662
rect 8898 -4718 8910 -4662
rect 8830 -4752 8910 -4718
rect 8830 -4808 8842 -4752
rect 8898 -4808 8910 -4752
rect 8830 -4820 8910 -4808
rect 220 -4972 390 -4960
rect 220 -5028 232 -4972
rect 288 -5028 322 -4972
rect 378 -5028 390 -4972
rect 220 -5040 390 -5028
rect 6300 -4972 6470 -4960
rect 6300 -5028 6312 -4972
rect 6368 -5028 6402 -4972
rect 6458 -5028 6470 -4972
rect 6300 -5040 6470 -5028
rect -110 -5082 60 -5070
rect -110 -5138 -98 -5082
rect -42 -5138 -8 -5082
rect 48 -5138 60 -5082
rect -110 -5150 60 -5138
rect -590 -5172 -490 -5150
rect -590 -5228 -568 -5172
rect -512 -5228 -490 -5172
rect -590 -5250 -490 -5228
<< via3 >>
rect 548 5158 612 5222
rect 668 5158 732 5222
rect 928 5158 992 5222
rect 1048 5158 1112 5222
rect 1308 5158 1372 5222
rect 1428 5158 1492 5222
rect 1688 5158 1752 5222
rect 1808 5158 1872 5222
rect 2068 5158 2132 5222
rect 2188 5158 2252 5222
rect 2448 5158 2512 5222
rect 2568 5158 2632 5222
rect 2828 5158 2892 5222
rect 2948 5158 3012 5222
rect 3208 5158 3272 5222
rect 3328 5158 3392 5222
rect 3588 5158 3652 5222
rect 3708 5158 3772 5222
rect 3968 5158 4032 5222
rect 4088 5158 4152 5222
rect 4728 5158 4792 5222
rect 4848 5158 4912 5222
rect 5108 5158 5172 5222
rect 5228 5158 5292 5222
rect 5488 5158 5552 5222
rect 5608 5158 5672 5222
rect 5868 5158 5932 5222
rect 5988 5158 6052 5222
rect 6248 5158 6312 5222
rect 6368 5158 6432 5222
rect 6628 5158 6692 5222
rect 6748 5158 6812 5222
rect 7008 5158 7072 5222
rect 7128 5158 7192 5222
rect 7388 5158 7452 5222
rect 7508 5158 7572 5222
rect 7768 5158 7832 5222
rect 7888 5158 7952 5222
rect 8148 5158 8212 5222
rect 8268 5158 8332 5222
<< metal4 >>
rect -590 5222 8910 5250
rect -590 5158 548 5222
rect 612 5158 668 5222
rect 732 5158 928 5222
rect 992 5158 1048 5222
rect 1112 5158 1308 5222
rect 1372 5158 1428 5222
rect 1492 5158 1688 5222
rect 1752 5158 1808 5222
rect 1872 5158 2068 5222
rect 2132 5158 2188 5222
rect 2252 5158 2448 5222
rect 2512 5158 2568 5222
rect 2632 5158 2828 5222
rect 2892 5158 2948 5222
rect 3012 5158 3208 5222
rect 3272 5158 3328 5222
rect 3392 5158 3588 5222
rect 3652 5158 3708 5222
rect 3772 5158 3968 5222
rect 4032 5158 4088 5222
rect 4152 5158 4728 5222
rect 4792 5158 4848 5222
rect 4912 5158 5108 5222
rect 5172 5158 5228 5222
rect 5292 5158 5488 5222
rect 5552 5158 5608 5222
rect 5672 5158 5868 5222
rect 5932 5158 5988 5222
rect 6052 5158 6248 5222
rect 6312 5158 6368 5222
rect 6432 5158 6628 5222
rect 6692 5158 6748 5222
rect 6812 5158 7008 5222
rect 7072 5158 7128 5222
rect 7192 5158 7388 5222
rect 7452 5158 7508 5222
rect 7572 5158 7768 5222
rect 7832 5158 7888 5222
rect 7952 5158 8148 5222
rect 8212 5158 8268 5222
rect 8332 5158 8910 5222
rect -590 5130 8910 5158
rect -590 -5050 -490 -4950
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_0
timestamp 1757161594
transform 0 1 1287 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_1
timestamp 1757161594
transform 0 1 147 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_2
timestamp 1757161594
transform 0 1 527 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_3
timestamp 1757161594
transform 0 1 907 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_4
timestamp 1757161594
transform 0 1 1667 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_5
timestamp 1757161594
transform 0 1 2047 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_6
timestamp 1757161594
transform 0 1 4327 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_7
timestamp 1757161594
transform 0 1 3947 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_8
timestamp 1757161594
transform 0 1 3567 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_9
timestamp 1757161594
transform 0 1 3187 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_10
timestamp 1757161594
transform 0 1 2807 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_11
timestamp 1757161594
transform 0 1 2427 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_12
timestamp 1757161594
transform 0 1 5847 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_13
timestamp 1757161594
transform 0 1 5087 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_14
timestamp 1757161594
transform 0 1 5467 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_15
timestamp 1757161594
transform 0 1 4707 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_16
timestamp 1757161594
transform 0 1 6227 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_17
timestamp 1757161594
transform 0 1 6607 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_18
timestamp 1757161594
transform 0 1 7367 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_19
timestamp 1757161594
transform 0 1 8507 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_20
timestamp 1757161594
transform 0 1 8127 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_21
timestamp 1757161594
transform 0 1 7747 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_22
timestamp 1757161594
transform 0 1 6987 1 0 -4572
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_23
timestamp 1757161594
transform 0 1 2047 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_24
timestamp 1757161594
transform 0 1 1287 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_25
timestamp 1757161594
transform 0 1 1667 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_26
timestamp 1757161594
transform 0 1 527 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_27
timestamp 1757161594
transform 0 1 907 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_28
timestamp 1757161594
transform 0 1 147 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_29
timestamp 1757161594
transform 0 1 4327 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_30
timestamp 1757161594
transform 0 1 3567 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_31
timestamp 1757161594
transform 0 1 3947 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_32
timestamp 1757161594
transform 0 1 2807 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_33
timestamp 1757161594
transform 0 1 3187 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_34
timestamp 1757161594
transform 0 1 2427 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_35
timestamp 1757161594
transform 0 1 6607 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_36
timestamp 1757161594
transform 0 1 5847 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_37
timestamp 1757161594
transform 0 1 6227 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_38
timestamp 1757161594
transform 0 1 5087 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_39
timestamp 1757161594
transform 0 1 5467 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_40
timestamp 1757161594
transform 0 1 4707 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_41
timestamp 1757161594
transform 0 1 8127 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_42
timestamp 1757161594
transform 0 1 8507 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_43
timestamp 1757161594
transform 0 1 7367 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_44
timestamp 1757161594
transform 0 1 7747 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_6WKBEZ  sky130_fd_pr__nfet_01v8_lvt_6WKBEZ_45
timestamp 1757161594
transform 0 1 6987 1 0 4528
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_0
timestamp 1757161594
transform 0 1 4327 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_1
timestamp 1757161594
transform 0 1 3567 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_2
timestamp 1757161594
transform 0 1 3947 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_3
timestamp 1757161594
transform 0 1 3187 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_4
timestamp 1757161594
transform 0 1 2807 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_5
timestamp 1757161594
transform 0 1 2427 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_6
timestamp 1757161594
transform 0 1 1287 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_7
timestamp 1757161594
transform 0 1 1667 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_8
timestamp 1757161594
transform 0 1 2047 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_9
timestamp 1757161594
transform 0 1 907 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_10
timestamp 1757161594
transform 0 1 527 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_12
timestamp 1757161594
transform 0 1 6987 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_13
timestamp 1757161594
transform 0 1 8127 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_14
timestamp 1757161594
transform 0 1 7747 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_15
timestamp 1757161594
transform 0 1 7367 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_16
timestamp 1757161594
transform 0 1 8507 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_17
timestamp 1757161594
transform 0 1 2047 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_18
timestamp 1757161594
transform 0 1 4707 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_19
timestamp 1757161594
transform 0 1 5087 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_20
timestamp 1757161594
transform 0 1 5467 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_21
timestamp 1757161594
transform 0 1 5847 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_22
timestamp 1757161594
transform 0 1 6227 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_23
timestamp 1757161594
transform 0 1 6607 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_24
timestamp 1757161594
transform 0 1 1667 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_25
timestamp 1757161594
transform 0 1 1287 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_26
timestamp 1757161594
transform 0 1 907 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_27
timestamp 1757161594
transform 0 1 527 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_29
timestamp 1757161594
transform 0 1 3947 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_30
timestamp 1757161594
transform 0 1 3567 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_31
timestamp 1757161594
transform 0 1 3187 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_32
timestamp 1757161594
transform 0 1 2807 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_33
timestamp 1757161594
transform 0 1 2427 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_34
timestamp 1757161594
transform 0 1 5847 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_35
timestamp 1757161594
transform 0 1 5467 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_36
timestamp 1757161594
transform 0 1 5087 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_37
timestamp 1757161594
transform 0 1 4707 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_38
timestamp 1757161594
transform 0 1 4327 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_39
timestamp 1757161594
transform 0 1 8127 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_40
timestamp 1757161594
transform 0 1 7747 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_41
timestamp 1757161594
transform 0 1 7367 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_42
timestamp 1757161594
transform 0 1 6987 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_43
timestamp 1757161594
transform 0 1 6607 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_44
timestamp 1757161594
transform 0 1 6227 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_45
timestamp 1757161594
transform 0 1 8507 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_46
timestamp 1757161594
transform 0 1 8507 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_47
timestamp 1757161594
transform 0 1 8127 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_48
timestamp 1757161594
transform 0 1 7747 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_49
timestamp 1757161594
transform 0 1 7367 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_50
timestamp 1757161594
transform 0 1 6987 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_51
timestamp 1757161594
transform 0 1 6607 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_52
timestamp 1757161594
transform 0 1 6227 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_53
timestamp 1757161594
transform 0 1 5847 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_54
timestamp 1757161594
transform 0 1 5467 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_55
timestamp 1757161594
transform 0 1 5087 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_56
timestamp 1757161594
transform 0 1 4707 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_57
timestamp 1757161594
transform 0 1 4327 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_58
timestamp 1757161594
transform 0 1 3947 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_59
timestamp 1757161594
transform 0 1 147 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_60
timestamp 1757161594
transform 0 1 147 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_61
timestamp 1757161594
transform 0 1 147 1 0 1068
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_62
timestamp 1757161594
transform 0 1 147 1 0 3248
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_63
timestamp 1757161594
transform 0 1 2047 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_64
timestamp 1757161594
transform 0 1 1667 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_65
timestamp 1757161594
transform 0 1 1287 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_66
timestamp 1757161594
transform 0 1 907 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_67
timestamp 1757161594
transform 0 1 2427 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_68
timestamp 1757161594
transform 0 1 527 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_69
timestamp 1757161594
transform 0 1 2047 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_70
timestamp 1757161594
transform 0 1 1667 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_71
timestamp 1757161594
transform 0 1 1287 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_72
timestamp 1757161594
transform 0 1 907 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_73
timestamp 1757161594
transform 0 1 527 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_75
timestamp 1757161594
transform 0 1 4327 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_76
timestamp 1757161594
transform 0 1 3947 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_77
timestamp 1757161594
transform 0 1 3567 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_78
timestamp 1757161594
transform 0 1 3187 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_79
timestamp 1757161594
transform 0 1 2807 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_80
timestamp 1757161594
transform 0 1 2427 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_81
timestamp 1757161594
transform 0 1 6607 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_82
timestamp 1757161594
transform 0 1 6227 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_83
timestamp 1757161594
transform 0 1 5847 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_84
timestamp 1757161594
transform 0 1 5467 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_85
timestamp 1757161594
transform 0 1 5087 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_86
timestamp 1757161594
transform 0 1 4707 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_87
timestamp 1757161594
transform 0 1 8507 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_88
timestamp 1757161594
transform 0 1 8127 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_89
timestamp 1757161594
transform 0 1 7747 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_90
timestamp 1757161594
transform 0 1 7367 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_91
timestamp 1757161594
transform 0 1 6987 1 0 -1112
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_93
timestamp 1757161594
transform 0 1 2807 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_94
timestamp 1757161594
transform 0 1 3187 1 0 -3292
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_lvt_F22EEM  sky130_fd_pr__nfet_01v8_lvt_F22EEM_95
timestamp 1757161594
transform 0 1 3567 1 0 -3292
box -1084 -157 1084 157
<< labels >>
flabel metal1 s 10 -5320 110 -5220 0 FreeSans 782 0 0 0 Vss
port 1 nsew
flabel metal1 s 10 5410 110 5510 0 FreeSans 782 0 0 0 Vss
port 1 nsew
flabel metal4 s -590 5130 -470 5250 0 FreeSans 782 0 0 0 Vbias2
port 2 nsew
<< end >>
