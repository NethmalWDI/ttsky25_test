magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -594 -198 594 164
<< pmoslvt >>
rect -500 -136 500 64
<< pdiff >>
rect -558 15 -500 64
rect -558 -19 -546 15
rect -512 -19 -500 15
rect -558 -53 -500 -19
rect -558 -87 -546 -53
rect -512 -87 -500 -53
rect -558 -136 -500 -87
rect 500 15 558 64
rect 500 -19 512 15
rect 546 -19 558 15
rect 500 -53 558 -19
rect 500 -87 512 -53
rect 546 -87 558 -53
rect 500 -136 558 -87
<< pdiffc >>
rect -546 -19 -512 15
rect -546 -87 -512 -53
rect 512 -19 546 15
rect 512 -87 546 -53
<< poly >>
rect -355 145 355 161
rect -355 128 -323 145
rect -500 111 -323 128
rect -289 111 -255 145
rect -221 111 -187 145
rect -153 111 -119 145
rect -85 111 -51 145
rect -17 111 17 145
rect 51 111 85 145
rect 119 111 153 145
rect 187 111 221 145
rect 255 111 289 145
rect 323 128 355 145
rect 323 111 500 128
rect -500 64 500 111
rect -500 -162 500 -136
<< polycont >>
rect -323 111 -289 145
rect -255 111 -221 145
rect -187 111 -153 145
rect -119 111 -85 145
rect -51 111 -17 145
rect 17 111 51 145
rect 85 111 119 145
rect 153 111 187 145
rect 221 111 255 145
rect 289 111 323 145
<< locali >>
rect -355 111 -323 145
rect -271 111 -255 145
rect -199 111 -187 145
rect -127 111 -119 145
rect -55 111 -51 145
rect 51 111 55 145
rect 119 111 127 145
rect 187 111 199 145
rect 255 111 271 145
rect 323 111 355 145
rect -546 17 -512 42
rect -546 -53 -512 -19
rect -546 -114 -512 -89
rect 512 17 546 42
rect 512 -53 546 -19
rect 512 -114 546 -89
<< viali >>
rect -305 111 -289 145
rect -289 111 -271 145
rect -233 111 -221 145
rect -221 111 -199 145
rect -161 111 -153 145
rect -153 111 -127 145
rect -89 111 -85 145
rect -85 111 -55 145
rect -17 111 17 145
rect 55 111 85 145
rect 85 111 89 145
rect 127 111 153 145
rect 153 111 161 145
rect 199 111 221 145
rect 221 111 233 145
rect 271 111 289 145
rect 289 111 305 145
rect -546 15 -512 17
rect -546 -17 -512 15
rect -546 -87 -512 -55
rect -546 -89 -512 -87
rect 512 15 546 17
rect 512 -17 546 15
rect 512 -87 546 -55
rect 512 -89 546 -87
<< metal1 >>
rect -351 145 351 151
rect -351 111 -305 145
rect -271 111 -233 145
rect -199 111 -161 145
rect -127 111 -89 145
rect -55 111 -17 145
rect 17 111 55 145
rect 89 111 127 145
rect 161 111 199 145
rect 233 111 271 145
rect 305 111 351 145
rect -351 105 351 111
rect -552 17 -506 38
rect -552 -17 -546 17
rect -512 -17 -506 17
rect -552 -55 -506 -17
rect -552 -89 -546 -55
rect -512 -89 -506 -55
rect -552 -110 -506 -89
rect 506 17 552 38
rect 506 -17 512 17
rect 546 -17 552 17
rect 506 -55 552 -17
rect 506 -89 512 -55
rect 546 -89 552 -55
rect 506 -110 552 -89
<< end >>
