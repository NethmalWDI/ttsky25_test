magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -396 -684 396 684
<< pmoslvt >>
rect -200 -536 200 464
<< pdiff >>
rect -258 423 -200 464
rect -258 389 -246 423
rect -212 389 -200 423
rect -258 355 -200 389
rect -258 321 -246 355
rect -212 321 -200 355
rect -258 287 -200 321
rect -258 253 -246 287
rect -212 253 -200 287
rect -258 219 -200 253
rect -258 185 -246 219
rect -212 185 -200 219
rect -258 151 -200 185
rect -258 117 -246 151
rect -212 117 -200 151
rect -258 83 -200 117
rect -258 49 -246 83
rect -212 49 -200 83
rect -258 15 -200 49
rect -258 -19 -246 15
rect -212 -19 -200 15
rect -258 -53 -200 -19
rect -258 -87 -246 -53
rect -212 -87 -200 -53
rect -258 -121 -200 -87
rect -258 -155 -246 -121
rect -212 -155 -200 -121
rect -258 -189 -200 -155
rect -258 -223 -246 -189
rect -212 -223 -200 -189
rect -258 -257 -200 -223
rect -258 -291 -246 -257
rect -212 -291 -200 -257
rect -258 -325 -200 -291
rect -258 -359 -246 -325
rect -212 -359 -200 -325
rect -258 -393 -200 -359
rect -258 -427 -246 -393
rect -212 -427 -200 -393
rect -258 -461 -200 -427
rect -258 -495 -246 -461
rect -212 -495 -200 -461
rect -258 -536 -200 -495
rect 200 423 258 464
rect 200 389 212 423
rect 246 389 258 423
rect 200 355 258 389
rect 200 321 212 355
rect 246 321 258 355
rect 200 287 258 321
rect 200 253 212 287
rect 246 253 258 287
rect 200 219 258 253
rect 200 185 212 219
rect 246 185 258 219
rect 200 151 258 185
rect 200 117 212 151
rect 246 117 258 151
rect 200 83 258 117
rect 200 49 212 83
rect 246 49 258 83
rect 200 15 258 49
rect 200 -19 212 15
rect 246 -19 258 15
rect 200 -53 258 -19
rect 200 -87 212 -53
rect 246 -87 258 -53
rect 200 -121 258 -87
rect 200 -155 212 -121
rect 246 -155 258 -121
rect 200 -189 258 -155
rect 200 -223 212 -189
rect 246 -223 258 -189
rect 200 -257 258 -223
rect 200 -291 212 -257
rect 246 -291 258 -257
rect 200 -325 258 -291
rect 200 -359 212 -325
rect 246 -359 258 -325
rect 200 -393 258 -359
rect 200 -427 212 -393
rect 246 -427 258 -393
rect 200 -461 258 -427
rect 200 -495 212 -461
rect 246 -495 258 -461
rect 200 -536 258 -495
<< pdiffc >>
rect -246 389 -212 423
rect -246 321 -212 355
rect -246 253 -212 287
rect -246 185 -212 219
rect -246 117 -212 151
rect -246 49 -212 83
rect -246 -19 -212 15
rect -246 -87 -212 -53
rect -246 -155 -212 -121
rect -246 -223 -212 -189
rect -246 -291 -212 -257
rect -246 -359 -212 -325
rect -246 -427 -212 -393
rect -246 -495 -212 -461
rect 212 389 246 423
rect 212 321 246 355
rect 212 253 246 287
rect 212 185 246 219
rect 212 117 246 151
rect 212 49 246 83
rect 212 -19 246 15
rect 212 -87 246 -53
rect 212 -155 246 -121
rect 212 -223 246 -189
rect 212 -291 246 -257
rect 212 -359 246 -325
rect 212 -427 246 -393
rect 212 -495 246 -461
<< nsubdiff >>
rect -360 614 360 648
rect -360 -614 -326 614
rect 326 -614 360 614
rect -360 -648 360 -614
<< poly >>
rect -200 545 200 561
rect -200 511 -153 545
rect -119 511 -85 545
rect -51 511 -17 545
rect 17 511 51 545
rect 85 511 119 545
rect 153 511 200 545
rect -200 464 200 511
rect -200 -562 200 -536
<< polycont >>
rect -153 511 -119 545
rect -85 511 -51 545
rect -17 511 17 545
rect 51 511 85 545
rect 119 511 153 545
<< locali >>
rect -360 614 360 648
rect -360 -614 -326 614
rect -200 511 -161 545
rect -119 511 -89 545
rect -51 511 -17 545
rect 17 511 51 545
rect 89 511 119 545
rect 161 511 200 545
rect -246 449 -212 468
rect -246 377 -212 389
rect -246 305 -212 321
rect -246 233 -212 253
rect -246 161 -212 185
rect -246 89 -212 117
rect -246 17 -212 49
rect -246 -53 -212 -19
rect -246 -121 -212 -89
rect -246 -189 -212 -161
rect -246 -257 -212 -233
rect -246 -325 -212 -305
rect -246 -393 -212 -377
rect -246 -461 -212 -449
rect -246 -540 -212 -521
rect 212 449 246 468
rect 212 377 246 389
rect 212 305 246 321
rect 212 233 246 253
rect 212 161 246 185
rect 212 89 246 117
rect 212 17 246 49
rect 212 -53 246 -19
rect 212 -121 246 -89
rect 212 -189 246 -161
rect 212 -257 246 -233
rect 212 -325 246 -305
rect 212 -393 246 -377
rect 212 -461 246 -449
rect 212 -540 246 -521
rect 326 -614 360 614
rect -360 -648 360 -614
<< viali >>
rect -161 511 -153 545
rect -153 511 -127 545
rect -89 511 -85 545
rect -85 511 -55 545
rect -17 511 17 545
rect 55 511 85 545
rect 85 511 89 545
rect 127 511 153 545
rect 153 511 161 545
rect -246 423 -212 449
rect -246 415 -212 423
rect -246 355 -212 377
rect -246 343 -212 355
rect -246 287 -212 305
rect -246 271 -212 287
rect -246 219 -212 233
rect -246 199 -212 219
rect -246 151 -212 161
rect -246 127 -212 151
rect -246 83 -212 89
rect -246 55 -212 83
rect -246 15 -212 17
rect -246 -17 -212 15
rect -246 -87 -212 -55
rect -246 -89 -212 -87
rect -246 -155 -212 -127
rect -246 -161 -212 -155
rect -246 -223 -212 -199
rect -246 -233 -212 -223
rect -246 -291 -212 -271
rect -246 -305 -212 -291
rect -246 -359 -212 -343
rect -246 -377 -212 -359
rect -246 -427 -212 -415
rect -246 -449 -212 -427
rect -246 -495 -212 -487
rect -246 -521 -212 -495
rect 212 423 246 449
rect 212 415 246 423
rect 212 355 246 377
rect 212 343 246 355
rect 212 287 246 305
rect 212 271 246 287
rect 212 219 246 233
rect 212 199 246 219
rect 212 151 246 161
rect 212 127 246 151
rect 212 83 246 89
rect 212 55 246 83
rect 212 15 246 17
rect 212 -17 246 15
rect 212 -87 246 -55
rect 212 -89 246 -87
rect 212 -155 246 -127
rect 212 -161 246 -155
rect 212 -223 246 -199
rect 212 -233 246 -223
rect 212 -291 246 -271
rect 212 -305 246 -291
rect 212 -359 246 -343
rect 212 -377 246 -359
rect 212 -427 246 -415
rect 212 -449 246 -427
rect 212 -495 246 -487
rect 212 -521 246 -495
<< metal1 >>
rect -196 545 196 551
rect -196 511 -161 545
rect -127 511 -89 545
rect -55 511 -17 545
rect 17 511 55 545
rect 89 511 127 545
rect 161 511 196 545
rect -196 505 196 511
rect -252 449 -206 464
rect -252 415 -246 449
rect -212 415 -206 449
rect -252 377 -206 415
rect -252 343 -246 377
rect -212 343 -206 377
rect -252 305 -206 343
rect -252 271 -246 305
rect -212 271 -206 305
rect -252 233 -206 271
rect -252 199 -246 233
rect -212 199 -206 233
rect -252 161 -206 199
rect -252 127 -246 161
rect -212 127 -206 161
rect -252 89 -206 127
rect -252 55 -246 89
rect -212 55 -206 89
rect -252 17 -206 55
rect -252 -17 -246 17
rect -212 -17 -206 17
rect -252 -55 -206 -17
rect -252 -89 -246 -55
rect -212 -89 -206 -55
rect -252 -127 -206 -89
rect -252 -161 -246 -127
rect -212 -161 -206 -127
rect -252 -199 -206 -161
rect -252 -233 -246 -199
rect -212 -233 -206 -199
rect -252 -271 -206 -233
rect -252 -305 -246 -271
rect -212 -305 -206 -271
rect -252 -343 -206 -305
rect -252 -377 -246 -343
rect -212 -377 -206 -343
rect -252 -415 -206 -377
rect -252 -449 -246 -415
rect -212 -449 -206 -415
rect -252 -487 -206 -449
rect -252 -521 -246 -487
rect -212 -521 -206 -487
rect -252 -536 -206 -521
rect 206 449 252 464
rect 206 415 212 449
rect 246 415 252 449
rect 206 377 252 415
rect 206 343 212 377
rect 246 343 252 377
rect 206 305 252 343
rect 206 271 212 305
rect 246 271 252 305
rect 206 233 252 271
rect 206 199 212 233
rect 246 199 252 233
rect 206 161 252 199
rect 206 127 212 161
rect 246 127 252 161
rect 206 89 252 127
rect 206 55 212 89
rect 246 55 252 89
rect 206 17 252 55
rect 206 -17 212 17
rect 246 -17 252 17
rect 206 -55 252 -17
rect 206 -89 212 -55
rect 246 -89 252 -55
rect 206 -127 252 -89
rect 206 -161 212 -127
rect 246 -161 252 -127
rect 206 -199 252 -161
rect 206 -233 212 -199
rect 246 -233 252 -199
rect 206 -271 252 -233
rect 206 -305 212 -271
rect 246 -305 252 -271
rect 206 -343 252 -305
rect 206 -377 212 -343
rect 246 -377 252 -343
rect 206 -415 252 -377
rect 206 -449 212 -415
rect 246 -449 252 -415
rect 206 -487 252 -449
rect 206 -521 212 -487
rect 246 -521 252 -487
rect 206 -536 252 -521
<< properties >>
string FIXED_BBOX -343 -631 343 631
<< end >>
