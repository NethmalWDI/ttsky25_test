magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< metal3 >>
rect -1186 512 1186 540
rect -1186 448 1102 512
rect 1166 448 1186 512
rect -1186 432 1186 448
rect -1186 368 1102 432
rect 1166 368 1186 432
rect -1186 352 1186 368
rect -1186 288 1102 352
rect 1166 288 1186 352
rect -1186 272 1186 288
rect -1186 208 1102 272
rect 1166 208 1186 272
rect -1186 192 1186 208
rect -1186 128 1102 192
rect 1166 128 1186 192
rect -1186 112 1186 128
rect -1186 48 1102 112
rect 1166 48 1186 112
rect -1186 32 1186 48
rect -1186 -32 1102 32
rect 1166 -32 1186 32
rect -1186 -48 1186 -32
rect -1186 -112 1102 -48
rect 1166 -112 1186 -48
rect -1186 -128 1186 -112
rect -1186 -192 1102 -128
rect 1166 -192 1186 -128
rect -1186 -208 1186 -192
rect -1186 -272 1102 -208
rect 1166 -272 1186 -208
rect -1186 -288 1186 -272
rect -1186 -352 1102 -288
rect 1166 -352 1186 -288
rect -1186 -368 1186 -352
rect -1186 -432 1102 -368
rect 1166 -432 1186 -368
rect -1186 -448 1186 -432
rect -1186 -512 1102 -448
rect 1166 -512 1186 -448
rect -1186 -540 1186 -512
<< via3 >>
rect 1102 448 1166 512
rect 1102 368 1166 432
rect 1102 288 1166 352
rect 1102 208 1166 272
rect 1102 128 1166 192
rect 1102 48 1166 112
rect 1102 -32 1166 32
rect 1102 -112 1166 -48
rect 1102 -192 1166 -128
rect 1102 -272 1166 -208
rect 1102 -352 1166 -288
rect 1102 -432 1166 -368
rect 1102 -512 1166 -448
<< mimcap >>
rect -1146 432 854 500
rect -1146 -432 -1098 432
rect 806 -432 854 432
rect -1146 -500 854 -432
<< mimcapcontact >>
rect -1098 -432 806 432
<< metal4 >>
rect 1086 512 1182 528
rect -1107 432 815 461
rect -1107 -432 -1098 432
rect 806 -432 815 432
rect -1107 -461 815 -432
rect 1086 448 1102 512
rect 1166 448 1182 512
rect 1086 432 1182 448
rect 1086 368 1102 432
rect 1166 368 1182 432
rect 1086 352 1182 368
rect 1086 288 1102 352
rect 1166 288 1182 352
rect 1086 272 1182 288
rect 1086 208 1102 272
rect 1166 208 1182 272
rect 1086 192 1182 208
rect 1086 128 1102 192
rect 1166 128 1182 192
rect 1086 112 1182 128
rect 1086 48 1102 112
rect 1166 48 1182 112
rect 1086 32 1182 48
rect 1086 -32 1102 32
rect 1166 -32 1182 32
rect 1086 -48 1182 -32
rect 1086 -112 1102 -48
rect 1166 -112 1182 -48
rect 1086 -128 1182 -112
rect 1086 -192 1102 -128
rect 1166 -192 1182 -128
rect 1086 -208 1182 -192
rect 1086 -272 1102 -208
rect 1166 -272 1182 -208
rect 1086 -288 1182 -272
rect 1086 -352 1102 -288
rect 1166 -352 1182 -288
rect 1086 -368 1182 -352
rect 1086 -432 1102 -368
rect 1166 -432 1182 -368
rect 1086 -448 1182 -432
rect 1086 -512 1102 -448
rect 1166 -512 1182 -448
rect 1086 -528 1182 -512
<< properties >>
string FIXED_BBOX -1186 -540 894 540
<< end >>
