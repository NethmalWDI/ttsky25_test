magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -153 -413 4063 9773
<< nsubdiff >>
rect -117 9703 -34 9737
rect 0 9703 34 9737
rect 68 9703 102 9737
rect 136 9703 170 9737
rect 204 9703 238 9737
rect 272 9703 306 9737
rect 340 9703 374 9737
rect 408 9703 442 9737
rect 476 9703 510 9737
rect 544 9703 578 9737
rect 612 9703 646 9737
rect 680 9703 714 9737
rect 748 9703 782 9737
rect 816 9703 850 9737
rect 884 9703 918 9737
rect 952 9703 986 9737
rect 1020 9703 1054 9737
rect 1088 9703 1122 9737
rect 1156 9703 1190 9737
rect 1224 9703 1258 9737
rect 1292 9703 1326 9737
rect 1360 9703 1394 9737
rect 1428 9703 1462 9737
rect 1496 9703 1530 9737
rect 1564 9703 1598 9737
rect 1632 9703 1666 9737
rect 1700 9703 1734 9737
rect 1768 9703 1802 9737
rect 1836 9703 1870 9737
rect 1904 9703 1938 9737
rect 1972 9703 2006 9737
rect 2040 9703 2074 9737
rect 2108 9703 2142 9737
rect 2176 9703 2210 9737
rect 2244 9703 2278 9737
rect 2312 9703 2346 9737
rect 2380 9703 2414 9737
rect 2448 9703 2482 9737
rect 2516 9703 2550 9737
rect 2584 9703 2618 9737
rect 2652 9703 2686 9737
rect 2720 9703 2754 9737
rect 2788 9703 2822 9737
rect 2856 9703 2890 9737
rect 2924 9703 2958 9737
rect 2992 9703 3026 9737
rect 3060 9703 3094 9737
rect 3128 9703 3162 9737
rect 3196 9703 3230 9737
rect 3264 9703 3298 9737
rect 3332 9703 3366 9737
rect 3400 9703 3434 9737
rect 3468 9703 3502 9737
rect 3536 9703 3570 9737
rect 3604 9703 3638 9737
rect 3672 9703 3706 9737
rect 3740 9703 3774 9737
rect 3808 9703 3842 9737
rect 3876 9703 3910 9737
rect 3944 9703 4027 9737
rect -117 9661 -83 9703
rect -117 9593 -83 9627
rect -117 9525 -83 9559
rect -117 9457 -83 9491
rect -117 9389 -83 9423
rect -117 9321 -83 9355
rect -117 9253 -83 9287
rect -117 9185 -83 9219
rect -117 9117 -83 9151
rect -117 9049 -83 9083
rect -117 8981 -83 9015
rect -117 8913 -83 8947
rect -117 8845 -83 8879
rect -117 8777 -83 8811
rect -117 8709 -83 8743
rect -117 8641 -83 8675
rect -117 8573 -83 8607
rect -117 8505 -83 8539
rect -117 8437 -83 8471
rect -117 8369 -83 8403
rect -117 8301 -83 8335
rect -117 8233 -83 8267
rect -117 8165 -83 8199
rect -117 8097 -83 8131
rect -117 8029 -83 8063
rect -117 7961 -83 7995
rect -117 7893 -83 7927
rect -117 7825 -83 7859
rect -117 7757 -83 7791
rect -117 7689 -83 7723
rect -117 7621 -83 7655
rect -117 7553 -83 7587
rect -117 7485 -83 7519
rect -117 7417 -83 7451
rect -117 7349 -83 7383
rect -117 7281 -83 7315
rect -117 7213 -83 7247
rect -117 7145 -83 7179
rect -117 7077 -83 7111
rect -117 7009 -83 7043
rect -117 6941 -83 6975
rect -117 6873 -83 6907
rect -117 6805 -83 6839
rect -117 6737 -83 6771
rect -117 6669 -83 6703
rect -117 6601 -83 6635
rect -117 6533 -83 6567
rect -117 6465 -83 6499
rect -117 6397 -83 6431
rect -117 6329 -83 6363
rect -117 6261 -83 6295
rect -117 6193 -83 6227
rect -117 6125 -83 6159
rect -117 6057 -83 6091
rect -117 5989 -83 6023
rect -117 5921 -83 5955
rect -117 5853 -83 5887
rect -117 5785 -83 5819
rect -117 5717 -83 5751
rect -117 5649 -83 5683
rect -117 5581 -83 5615
rect -117 5513 -83 5547
rect -117 5445 -83 5479
rect -117 5377 -83 5411
rect -117 5309 -83 5343
rect -117 5241 -83 5275
rect -117 5173 -83 5207
rect -117 5105 -83 5139
rect -117 5037 -83 5071
rect -117 4969 -83 5003
rect -117 4901 -83 4935
rect -117 4833 -83 4867
rect -117 4765 -83 4799
rect -117 4697 -83 4731
rect -117 4629 -83 4663
rect -117 4561 -83 4595
rect -117 4493 -83 4527
rect -117 4425 -83 4459
rect -117 4357 -83 4391
rect -117 4289 -83 4323
rect -117 4221 -83 4255
rect -117 4153 -83 4187
rect -117 4085 -83 4119
rect -117 4017 -83 4051
rect -117 3949 -83 3983
rect -117 3881 -83 3915
rect -117 3813 -83 3847
rect -117 3745 -83 3779
rect -117 3677 -83 3711
rect -117 3609 -83 3643
rect -117 3541 -83 3575
rect -117 3473 -83 3507
rect -117 3405 -83 3439
rect -117 3337 -83 3371
rect -117 3269 -83 3303
rect -117 3201 -83 3235
rect -117 3133 -83 3167
rect -117 3065 -83 3099
rect -117 2997 -83 3031
rect -117 2929 -83 2963
rect -117 2861 -83 2895
rect -117 2793 -83 2827
rect -117 2725 -83 2759
rect -117 2657 -83 2691
rect -117 2589 -83 2623
rect -117 2521 -83 2555
rect -117 2453 -83 2487
rect -117 2385 -83 2419
rect -117 2317 -83 2351
rect -117 2249 -83 2283
rect -117 2181 -83 2215
rect -117 2113 -83 2147
rect -117 2045 -83 2079
rect -117 1977 -83 2011
rect -117 1909 -83 1943
rect -117 1841 -83 1875
rect -117 1773 -83 1807
rect -117 1705 -83 1739
rect -117 1637 -83 1671
rect -117 1569 -83 1603
rect -117 1501 -83 1535
rect -117 1433 -83 1467
rect -117 1365 -83 1399
rect -117 1297 -83 1331
rect -117 1229 -83 1263
rect -117 1161 -83 1195
rect -117 1093 -83 1127
rect -117 1025 -83 1059
rect -117 957 -83 991
rect -117 889 -83 923
rect -117 821 -83 855
rect -117 753 -83 787
rect -117 685 -83 719
rect -117 617 -83 651
rect -117 549 -83 583
rect -117 481 -83 515
rect -117 413 -83 447
rect -117 345 -83 379
rect -117 277 -83 311
rect -117 209 -83 243
rect -117 141 -83 175
rect -117 73 -83 107
rect -117 5 -83 39
rect -117 -63 -83 -29
rect -117 -131 -83 -97
rect -117 -199 -83 -165
rect -117 -267 -83 -233
rect -117 -343 -83 -301
rect 3993 9661 4027 9703
rect 3993 9593 4027 9627
rect 3993 9525 4027 9559
rect 3993 9457 4027 9491
rect 3993 9389 4027 9423
rect 3993 9321 4027 9355
rect 3993 9253 4027 9287
rect 3993 9185 4027 9219
rect 3993 9117 4027 9151
rect 3993 9049 4027 9083
rect 3993 8981 4027 9015
rect 3993 8913 4027 8947
rect 3993 8845 4027 8879
rect 3993 8777 4027 8811
rect 3993 8709 4027 8743
rect 3993 8641 4027 8675
rect 3993 8573 4027 8607
rect 3993 8505 4027 8539
rect 3993 8437 4027 8471
rect 3993 8369 4027 8403
rect 3993 8301 4027 8335
rect 3993 8233 4027 8267
rect 3993 8165 4027 8199
rect 3993 8097 4027 8131
rect 3993 8029 4027 8063
rect 3993 7961 4027 7995
rect 3993 7893 4027 7927
rect 3993 7825 4027 7859
rect 3993 7757 4027 7791
rect 3993 7689 4027 7723
rect 3993 7621 4027 7655
rect 3993 7553 4027 7587
rect 3993 7485 4027 7519
rect 3993 7417 4027 7451
rect 3993 7349 4027 7383
rect 3993 7281 4027 7315
rect 3993 7213 4027 7247
rect 3993 7145 4027 7179
rect 3993 7077 4027 7111
rect 3993 7009 4027 7043
rect 3993 6941 4027 6975
rect 3993 6873 4027 6907
rect 3993 6805 4027 6839
rect 3993 6737 4027 6771
rect 3993 6669 4027 6703
rect 3993 6601 4027 6635
rect 3993 6533 4027 6567
rect 3993 6465 4027 6499
rect 3993 6397 4027 6431
rect 3993 6329 4027 6363
rect 3993 6261 4027 6295
rect 3993 6193 4027 6227
rect 3993 6125 4027 6159
rect 3993 6057 4027 6091
rect 3993 5989 4027 6023
rect 3993 5921 4027 5955
rect 3993 5853 4027 5887
rect 3993 5785 4027 5819
rect 3993 5717 4027 5751
rect 3993 5649 4027 5683
rect 3993 5581 4027 5615
rect 3993 5513 4027 5547
rect 3993 5445 4027 5479
rect 3993 5377 4027 5411
rect 3993 5309 4027 5343
rect 3993 5241 4027 5275
rect 3993 5173 4027 5207
rect 3993 5105 4027 5139
rect 3993 5037 4027 5071
rect 3993 4969 4027 5003
rect 3993 4901 4027 4935
rect 3993 4833 4027 4867
rect 3993 4765 4027 4799
rect 3993 4697 4027 4731
rect 3993 4629 4027 4663
rect 3993 4561 4027 4595
rect 3993 4493 4027 4527
rect 3993 4425 4027 4459
rect 3993 4357 4027 4391
rect 3993 4289 4027 4323
rect 3993 4221 4027 4255
rect 3993 4153 4027 4187
rect 3993 4085 4027 4119
rect 3993 4017 4027 4051
rect 3993 3949 4027 3983
rect 3993 3881 4027 3915
rect 3993 3813 4027 3847
rect 3993 3745 4027 3779
rect 3993 3677 4027 3711
rect 3993 3609 4027 3643
rect 3993 3541 4027 3575
rect 3993 3473 4027 3507
rect 3993 3405 4027 3439
rect 3993 3337 4027 3371
rect 3993 3269 4027 3303
rect 3993 3201 4027 3235
rect 3993 3133 4027 3167
rect 3993 3065 4027 3099
rect 3993 2997 4027 3031
rect 3993 2929 4027 2963
rect 3993 2861 4027 2895
rect 3993 2793 4027 2827
rect 3993 2725 4027 2759
rect 3993 2657 4027 2691
rect 3993 2589 4027 2623
rect 3993 2521 4027 2555
rect 3993 2453 4027 2487
rect 3993 2385 4027 2419
rect 3993 2317 4027 2351
rect 3993 2249 4027 2283
rect 3993 2181 4027 2215
rect 3993 2113 4027 2147
rect 3993 2045 4027 2079
rect 3993 1977 4027 2011
rect 3993 1909 4027 1943
rect 3993 1841 4027 1875
rect 3993 1773 4027 1807
rect 3993 1705 4027 1739
rect 3993 1637 4027 1671
rect 3993 1569 4027 1603
rect 3993 1501 4027 1535
rect 3993 1433 4027 1467
rect 3993 1365 4027 1399
rect 3993 1297 4027 1331
rect 3993 1229 4027 1263
rect 3993 1161 4027 1195
rect 3993 1093 4027 1127
rect 3993 1025 4027 1059
rect 3993 957 4027 991
rect 3993 889 4027 923
rect 3993 821 4027 855
rect 3993 753 4027 787
rect 3993 685 4027 719
rect 3993 617 4027 651
rect 3993 549 4027 583
rect 3993 481 4027 515
rect 3993 413 4027 447
rect 3993 345 4027 379
rect 3993 277 4027 311
rect 3993 209 4027 243
rect 3993 141 4027 175
rect 3993 73 4027 107
rect 3993 5 4027 39
rect 3993 -63 4027 -29
rect 3993 -131 4027 -97
rect 3993 -199 4027 -165
rect 3993 -267 4027 -233
rect 3993 -343 4027 -301
rect -117 -377 -34 -343
rect 0 -377 34 -343
rect 68 -377 102 -343
rect 136 -377 170 -343
rect 204 -377 238 -343
rect 272 -377 306 -343
rect 340 -377 374 -343
rect 408 -377 442 -343
rect 476 -377 510 -343
rect 544 -377 578 -343
rect 612 -377 646 -343
rect 680 -377 714 -343
rect 748 -377 782 -343
rect 816 -377 850 -343
rect 884 -377 918 -343
rect 952 -377 986 -343
rect 1020 -377 1054 -343
rect 1088 -377 1122 -343
rect 1156 -377 1190 -343
rect 1224 -377 1258 -343
rect 1292 -377 1326 -343
rect 1360 -377 1394 -343
rect 1428 -377 1462 -343
rect 1496 -377 1530 -343
rect 1564 -377 1598 -343
rect 1632 -377 1666 -343
rect 1700 -377 1734 -343
rect 1768 -377 1802 -343
rect 1836 -377 1870 -343
rect 1904 -377 1938 -343
rect 1972 -377 2006 -343
rect 2040 -377 2074 -343
rect 2108 -377 2142 -343
rect 2176 -377 2210 -343
rect 2244 -377 2278 -343
rect 2312 -377 2346 -343
rect 2380 -377 2414 -343
rect 2448 -377 2482 -343
rect 2516 -377 2550 -343
rect 2584 -377 2618 -343
rect 2652 -377 2686 -343
rect 2720 -377 2754 -343
rect 2788 -377 2822 -343
rect 2856 -377 2890 -343
rect 2924 -377 2958 -343
rect 2992 -377 3026 -343
rect 3060 -377 3094 -343
rect 3128 -377 3162 -343
rect 3196 -377 3230 -343
rect 3264 -377 3298 -343
rect 3332 -377 3366 -343
rect 3400 -377 3434 -343
rect 3468 -377 3502 -343
rect 3536 -377 3570 -343
rect 3604 -377 3638 -343
rect 3672 -377 3706 -343
rect 3740 -377 3774 -343
rect 3808 -377 3842 -343
rect 3876 -377 3910 -343
rect 3944 -377 4027 -343
<< nsubdiffcont >>
rect -34 9703 0 9737
rect 34 9703 68 9737
rect 102 9703 136 9737
rect 170 9703 204 9737
rect 238 9703 272 9737
rect 306 9703 340 9737
rect 374 9703 408 9737
rect 442 9703 476 9737
rect 510 9703 544 9737
rect 578 9703 612 9737
rect 646 9703 680 9737
rect 714 9703 748 9737
rect 782 9703 816 9737
rect 850 9703 884 9737
rect 918 9703 952 9737
rect 986 9703 1020 9737
rect 1054 9703 1088 9737
rect 1122 9703 1156 9737
rect 1190 9703 1224 9737
rect 1258 9703 1292 9737
rect 1326 9703 1360 9737
rect 1394 9703 1428 9737
rect 1462 9703 1496 9737
rect 1530 9703 1564 9737
rect 1598 9703 1632 9737
rect 1666 9703 1700 9737
rect 1734 9703 1768 9737
rect 1802 9703 1836 9737
rect 1870 9703 1904 9737
rect 1938 9703 1972 9737
rect 2006 9703 2040 9737
rect 2074 9703 2108 9737
rect 2142 9703 2176 9737
rect 2210 9703 2244 9737
rect 2278 9703 2312 9737
rect 2346 9703 2380 9737
rect 2414 9703 2448 9737
rect 2482 9703 2516 9737
rect 2550 9703 2584 9737
rect 2618 9703 2652 9737
rect 2686 9703 2720 9737
rect 2754 9703 2788 9737
rect 2822 9703 2856 9737
rect 2890 9703 2924 9737
rect 2958 9703 2992 9737
rect 3026 9703 3060 9737
rect 3094 9703 3128 9737
rect 3162 9703 3196 9737
rect 3230 9703 3264 9737
rect 3298 9703 3332 9737
rect 3366 9703 3400 9737
rect 3434 9703 3468 9737
rect 3502 9703 3536 9737
rect 3570 9703 3604 9737
rect 3638 9703 3672 9737
rect 3706 9703 3740 9737
rect 3774 9703 3808 9737
rect 3842 9703 3876 9737
rect 3910 9703 3944 9737
rect -117 9627 -83 9661
rect -117 9559 -83 9593
rect -117 9491 -83 9525
rect -117 9423 -83 9457
rect -117 9355 -83 9389
rect -117 9287 -83 9321
rect -117 9219 -83 9253
rect -117 9151 -83 9185
rect -117 9083 -83 9117
rect -117 9015 -83 9049
rect -117 8947 -83 8981
rect -117 8879 -83 8913
rect -117 8811 -83 8845
rect -117 8743 -83 8777
rect -117 8675 -83 8709
rect -117 8607 -83 8641
rect -117 8539 -83 8573
rect -117 8471 -83 8505
rect -117 8403 -83 8437
rect -117 8335 -83 8369
rect -117 8267 -83 8301
rect -117 8199 -83 8233
rect -117 8131 -83 8165
rect -117 8063 -83 8097
rect -117 7995 -83 8029
rect -117 7927 -83 7961
rect -117 7859 -83 7893
rect -117 7791 -83 7825
rect -117 7723 -83 7757
rect -117 7655 -83 7689
rect -117 7587 -83 7621
rect -117 7519 -83 7553
rect -117 7451 -83 7485
rect -117 7383 -83 7417
rect -117 7315 -83 7349
rect -117 7247 -83 7281
rect -117 7179 -83 7213
rect -117 7111 -83 7145
rect -117 7043 -83 7077
rect -117 6975 -83 7009
rect -117 6907 -83 6941
rect -117 6839 -83 6873
rect -117 6771 -83 6805
rect -117 6703 -83 6737
rect -117 6635 -83 6669
rect -117 6567 -83 6601
rect -117 6499 -83 6533
rect -117 6431 -83 6465
rect -117 6363 -83 6397
rect -117 6295 -83 6329
rect -117 6227 -83 6261
rect -117 6159 -83 6193
rect -117 6091 -83 6125
rect -117 6023 -83 6057
rect -117 5955 -83 5989
rect -117 5887 -83 5921
rect -117 5819 -83 5853
rect -117 5751 -83 5785
rect -117 5683 -83 5717
rect -117 5615 -83 5649
rect -117 5547 -83 5581
rect -117 5479 -83 5513
rect -117 5411 -83 5445
rect -117 5343 -83 5377
rect -117 5275 -83 5309
rect -117 5207 -83 5241
rect -117 5139 -83 5173
rect -117 5071 -83 5105
rect -117 5003 -83 5037
rect -117 4935 -83 4969
rect -117 4867 -83 4901
rect -117 4799 -83 4833
rect -117 4731 -83 4765
rect -117 4663 -83 4697
rect -117 4595 -83 4629
rect -117 4527 -83 4561
rect -117 4459 -83 4493
rect -117 4391 -83 4425
rect -117 4323 -83 4357
rect -117 4255 -83 4289
rect -117 4187 -83 4221
rect -117 4119 -83 4153
rect -117 4051 -83 4085
rect -117 3983 -83 4017
rect -117 3915 -83 3949
rect -117 3847 -83 3881
rect -117 3779 -83 3813
rect -117 3711 -83 3745
rect -117 3643 -83 3677
rect -117 3575 -83 3609
rect -117 3507 -83 3541
rect -117 3439 -83 3473
rect -117 3371 -83 3405
rect -117 3303 -83 3337
rect -117 3235 -83 3269
rect -117 3167 -83 3201
rect -117 3099 -83 3133
rect -117 3031 -83 3065
rect -117 2963 -83 2997
rect -117 2895 -83 2929
rect -117 2827 -83 2861
rect -117 2759 -83 2793
rect -117 2691 -83 2725
rect -117 2623 -83 2657
rect -117 2555 -83 2589
rect -117 2487 -83 2521
rect -117 2419 -83 2453
rect -117 2351 -83 2385
rect -117 2283 -83 2317
rect -117 2215 -83 2249
rect -117 2147 -83 2181
rect -117 2079 -83 2113
rect -117 2011 -83 2045
rect -117 1943 -83 1977
rect -117 1875 -83 1909
rect -117 1807 -83 1841
rect -117 1739 -83 1773
rect -117 1671 -83 1705
rect -117 1603 -83 1637
rect -117 1535 -83 1569
rect -117 1467 -83 1501
rect -117 1399 -83 1433
rect -117 1331 -83 1365
rect -117 1263 -83 1297
rect -117 1195 -83 1229
rect -117 1127 -83 1161
rect -117 1059 -83 1093
rect -117 991 -83 1025
rect -117 923 -83 957
rect -117 855 -83 889
rect -117 787 -83 821
rect -117 719 -83 753
rect -117 651 -83 685
rect -117 583 -83 617
rect -117 515 -83 549
rect -117 447 -83 481
rect -117 379 -83 413
rect -117 311 -83 345
rect -117 243 -83 277
rect -117 175 -83 209
rect -117 107 -83 141
rect -117 39 -83 73
rect -117 -29 -83 5
rect -117 -97 -83 -63
rect -117 -165 -83 -131
rect -117 -233 -83 -199
rect -117 -301 -83 -267
rect 3993 9627 4027 9661
rect 3993 9559 4027 9593
rect 3993 9491 4027 9525
rect 3993 9423 4027 9457
rect 3993 9355 4027 9389
rect 3993 9287 4027 9321
rect 3993 9219 4027 9253
rect 3993 9151 4027 9185
rect 3993 9083 4027 9117
rect 3993 9015 4027 9049
rect 3993 8947 4027 8981
rect 3993 8879 4027 8913
rect 3993 8811 4027 8845
rect 3993 8743 4027 8777
rect 3993 8675 4027 8709
rect 3993 8607 4027 8641
rect 3993 8539 4027 8573
rect 3993 8471 4027 8505
rect 3993 8403 4027 8437
rect 3993 8335 4027 8369
rect 3993 8267 4027 8301
rect 3993 8199 4027 8233
rect 3993 8131 4027 8165
rect 3993 8063 4027 8097
rect 3993 7995 4027 8029
rect 3993 7927 4027 7961
rect 3993 7859 4027 7893
rect 3993 7791 4027 7825
rect 3993 7723 4027 7757
rect 3993 7655 4027 7689
rect 3993 7587 4027 7621
rect 3993 7519 4027 7553
rect 3993 7451 4027 7485
rect 3993 7383 4027 7417
rect 3993 7315 4027 7349
rect 3993 7247 4027 7281
rect 3993 7179 4027 7213
rect 3993 7111 4027 7145
rect 3993 7043 4027 7077
rect 3993 6975 4027 7009
rect 3993 6907 4027 6941
rect 3993 6839 4027 6873
rect 3993 6771 4027 6805
rect 3993 6703 4027 6737
rect 3993 6635 4027 6669
rect 3993 6567 4027 6601
rect 3993 6499 4027 6533
rect 3993 6431 4027 6465
rect 3993 6363 4027 6397
rect 3993 6295 4027 6329
rect 3993 6227 4027 6261
rect 3993 6159 4027 6193
rect 3993 6091 4027 6125
rect 3993 6023 4027 6057
rect 3993 5955 4027 5989
rect 3993 5887 4027 5921
rect 3993 5819 4027 5853
rect 3993 5751 4027 5785
rect 3993 5683 4027 5717
rect 3993 5615 4027 5649
rect 3993 5547 4027 5581
rect 3993 5479 4027 5513
rect 3993 5411 4027 5445
rect 3993 5343 4027 5377
rect 3993 5275 4027 5309
rect 3993 5207 4027 5241
rect 3993 5139 4027 5173
rect 3993 5071 4027 5105
rect 3993 5003 4027 5037
rect 3993 4935 4027 4969
rect 3993 4867 4027 4901
rect 3993 4799 4027 4833
rect 3993 4731 4027 4765
rect 3993 4663 4027 4697
rect 3993 4595 4027 4629
rect 3993 4527 4027 4561
rect 3993 4459 4027 4493
rect 3993 4391 4027 4425
rect 3993 4323 4027 4357
rect 3993 4255 4027 4289
rect 3993 4187 4027 4221
rect 3993 4119 4027 4153
rect 3993 4051 4027 4085
rect 3993 3983 4027 4017
rect 3993 3915 4027 3949
rect 3993 3847 4027 3881
rect 3993 3779 4027 3813
rect 3993 3711 4027 3745
rect 3993 3643 4027 3677
rect 3993 3575 4027 3609
rect 3993 3507 4027 3541
rect 3993 3439 4027 3473
rect 3993 3371 4027 3405
rect 3993 3303 4027 3337
rect 3993 3235 4027 3269
rect 3993 3167 4027 3201
rect 3993 3099 4027 3133
rect 3993 3031 4027 3065
rect 3993 2963 4027 2997
rect 3993 2895 4027 2929
rect 3993 2827 4027 2861
rect 3993 2759 4027 2793
rect 3993 2691 4027 2725
rect 3993 2623 4027 2657
rect 3993 2555 4027 2589
rect 3993 2487 4027 2521
rect 3993 2419 4027 2453
rect 3993 2351 4027 2385
rect 3993 2283 4027 2317
rect 3993 2215 4027 2249
rect 3993 2147 4027 2181
rect 3993 2079 4027 2113
rect 3993 2011 4027 2045
rect 3993 1943 4027 1977
rect 3993 1875 4027 1909
rect 3993 1807 4027 1841
rect 3993 1739 4027 1773
rect 3993 1671 4027 1705
rect 3993 1603 4027 1637
rect 3993 1535 4027 1569
rect 3993 1467 4027 1501
rect 3993 1399 4027 1433
rect 3993 1331 4027 1365
rect 3993 1263 4027 1297
rect 3993 1195 4027 1229
rect 3993 1127 4027 1161
rect 3993 1059 4027 1093
rect 3993 991 4027 1025
rect 3993 923 4027 957
rect 3993 855 4027 889
rect 3993 787 4027 821
rect 3993 719 4027 753
rect 3993 651 4027 685
rect 3993 583 4027 617
rect 3993 515 4027 549
rect 3993 447 4027 481
rect 3993 379 4027 413
rect 3993 311 4027 345
rect 3993 243 4027 277
rect 3993 175 4027 209
rect 3993 107 4027 141
rect 3993 39 4027 73
rect 3993 -29 4027 5
rect 3993 -97 4027 -63
rect 3993 -165 4027 -131
rect 3993 -233 4027 -199
rect 3993 -301 4027 -267
rect -34 -377 0 -343
rect 34 -377 68 -343
rect 102 -377 136 -343
rect 170 -377 204 -343
rect 238 -377 272 -343
rect 306 -377 340 -343
rect 374 -377 408 -343
rect 442 -377 476 -343
rect 510 -377 544 -343
rect 578 -377 612 -343
rect 646 -377 680 -343
rect 714 -377 748 -343
rect 782 -377 816 -343
rect 850 -377 884 -343
rect 918 -377 952 -343
rect 986 -377 1020 -343
rect 1054 -377 1088 -343
rect 1122 -377 1156 -343
rect 1190 -377 1224 -343
rect 1258 -377 1292 -343
rect 1326 -377 1360 -343
rect 1394 -377 1428 -343
rect 1462 -377 1496 -343
rect 1530 -377 1564 -343
rect 1598 -377 1632 -343
rect 1666 -377 1700 -343
rect 1734 -377 1768 -343
rect 1802 -377 1836 -343
rect 1870 -377 1904 -343
rect 1938 -377 1972 -343
rect 2006 -377 2040 -343
rect 2074 -377 2108 -343
rect 2142 -377 2176 -343
rect 2210 -377 2244 -343
rect 2278 -377 2312 -343
rect 2346 -377 2380 -343
rect 2414 -377 2448 -343
rect 2482 -377 2516 -343
rect 2550 -377 2584 -343
rect 2618 -377 2652 -343
rect 2686 -377 2720 -343
rect 2754 -377 2788 -343
rect 2822 -377 2856 -343
rect 2890 -377 2924 -343
rect 2958 -377 2992 -343
rect 3026 -377 3060 -343
rect 3094 -377 3128 -343
rect 3162 -377 3196 -343
rect 3230 -377 3264 -343
rect 3298 -377 3332 -343
rect 3366 -377 3400 -343
rect 3434 -377 3468 -343
rect 3502 -377 3536 -343
rect 3570 -377 3604 -343
rect 3638 -377 3672 -343
rect 3706 -377 3740 -343
rect 3774 -377 3808 -343
rect 3842 -377 3876 -343
rect 3910 -377 3944 -343
<< locali >>
rect -117 9703 -34 9737
rect 0 9703 34 9737
rect 68 9703 102 9737
rect 136 9703 170 9737
rect 204 9703 238 9737
rect 272 9703 306 9737
rect 340 9703 374 9737
rect 408 9703 442 9737
rect 476 9703 510 9737
rect 544 9703 578 9737
rect 612 9703 646 9737
rect 680 9703 714 9737
rect 748 9703 782 9737
rect 816 9703 850 9737
rect 884 9703 918 9737
rect 952 9703 986 9737
rect 1020 9703 1054 9737
rect 1088 9703 1122 9737
rect 1156 9703 1190 9737
rect 1224 9703 1258 9737
rect 1292 9703 1326 9737
rect 1360 9703 1394 9737
rect 1428 9703 1462 9737
rect 1496 9703 1530 9737
rect 1564 9703 1598 9737
rect 1632 9703 1666 9737
rect 1700 9703 1734 9737
rect 1768 9703 1802 9737
rect 1836 9703 1870 9737
rect 1904 9703 1938 9737
rect 1972 9703 2006 9737
rect 2040 9703 2074 9737
rect 2108 9703 2142 9737
rect 2176 9703 2210 9737
rect 2244 9703 2278 9737
rect 2312 9703 2346 9737
rect 2380 9703 2414 9737
rect 2448 9703 2482 9737
rect 2516 9703 2550 9737
rect 2584 9703 2618 9737
rect 2652 9703 2686 9737
rect 2720 9703 2754 9737
rect 2788 9703 2822 9737
rect 2856 9703 2890 9737
rect 2924 9703 2958 9737
rect 2992 9703 3026 9737
rect 3060 9703 3094 9737
rect 3128 9703 3162 9737
rect 3196 9703 3230 9737
rect 3264 9703 3298 9737
rect 3332 9703 3366 9737
rect 3400 9703 3434 9737
rect 3468 9703 3502 9737
rect 3536 9703 3570 9737
rect 3604 9703 3638 9737
rect 3672 9703 3706 9737
rect 3740 9703 3774 9737
rect 3808 9703 3842 9737
rect 3876 9703 3910 9737
rect 3944 9703 4027 9737
rect -117 9661 -83 9703
rect -117 9593 -83 9627
rect -117 9525 -83 9559
rect -117 9457 -83 9491
rect -117 9389 -83 9423
rect -117 9321 -83 9355
rect -117 9253 -83 9287
rect -117 9185 -83 9219
rect -117 9117 -83 9151
rect -117 9049 -83 9083
rect -117 8981 -83 9015
rect -117 8913 -83 8947
rect -117 8845 -83 8879
rect -117 8777 -83 8811
rect -117 8709 -83 8743
rect -117 8641 -83 8675
rect -117 8573 -83 8607
rect -117 8505 -83 8539
rect -117 8437 -83 8471
rect -117 8369 -83 8403
rect -117 8301 -83 8335
rect -117 8233 -83 8267
rect -117 8165 -83 8199
rect -117 8097 -83 8131
rect -117 8029 -83 8063
rect -117 7961 -83 7995
rect -117 7893 -83 7927
rect -117 7825 -83 7859
rect -117 7757 -83 7791
rect -117 7689 -83 7723
rect -117 7621 -83 7655
rect -117 7553 -83 7587
rect -117 7485 -83 7519
rect -117 7417 -83 7451
rect -117 7349 -83 7383
rect -117 7281 -83 7315
rect -117 7213 -83 7247
rect -117 7145 -83 7179
rect -117 7077 -83 7111
rect -117 7009 -83 7043
rect -117 6941 -83 6975
rect -117 6873 -83 6907
rect -117 6805 -83 6839
rect -117 6737 -83 6771
rect -117 6669 -83 6703
rect -117 6601 -83 6635
rect -117 6533 -83 6567
rect -117 6465 -83 6499
rect -117 6397 -83 6431
rect -117 6329 -83 6363
rect -117 6261 -83 6295
rect -117 6193 -83 6227
rect -117 6125 -83 6159
rect -117 6057 -83 6091
rect -117 5989 -83 6023
rect -117 5921 -83 5955
rect -117 5853 -83 5887
rect -117 5785 -83 5819
rect -117 5717 -83 5751
rect -117 5649 -83 5683
rect -117 5581 -83 5615
rect -117 5513 -83 5547
rect -117 5445 -83 5479
rect -117 5377 -83 5411
rect -117 5309 -83 5343
rect -117 5241 -83 5275
rect -117 5173 -83 5207
rect -117 5105 -83 5139
rect -117 5037 -83 5071
rect -117 4969 -83 5003
rect -117 4901 -83 4935
rect -117 4833 -83 4867
rect -117 4765 -83 4799
rect -117 4697 -83 4731
rect -117 4629 -83 4663
rect -117 4561 -83 4595
rect -117 4493 -83 4527
rect -117 4425 -83 4459
rect -117 4357 -83 4391
rect -117 4289 -83 4323
rect -117 4221 -83 4255
rect -117 4153 -83 4187
rect -117 4085 -83 4119
rect -117 4017 -83 4051
rect -117 3949 -83 3983
rect -117 3881 -83 3915
rect -117 3813 -83 3847
rect -117 3745 -83 3779
rect -117 3677 -83 3711
rect -117 3609 -83 3643
rect -117 3541 -83 3575
rect -117 3473 -83 3507
rect -117 3405 -83 3439
rect -117 3337 -83 3371
rect -117 3269 -83 3303
rect -117 3201 -83 3235
rect -117 3133 -83 3167
rect -117 3065 -83 3099
rect -117 2997 -83 3031
rect -117 2929 -83 2963
rect -117 2861 -83 2895
rect -117 2793 -83 2827
rect -117 2725 -83 2759
rect -117 2657 -83 2691
rect -117 2589 -83 2623
rect -117 2521 -83 2555
rect -117 2453 -83 2487
rect -117 2385 -83 2419
rect -117 2317 -83 2351
rect -117 2249 -83 2283
rect -117 2181 -83 2215
rect -117 2113 -83 2147
rect -117 2045 -83 2079
rect -117 1977 -83 2011
rect -117 1909 -83 1943
rect -117 1841 -83 1875
rect -117 1773 -83 1807
rect -117 1705 -83 1739
rect -117 1637 -83 1671
rect -117 1569 -83 1603
rect -117 1501 -83 1535
rect -117 1433 -83 1467
rect -117 1365 -83 1399
rect -117 1297 -83 1331
rect -117 1229 -83 1263
rect -117 1161 -83 1195
rect -117 1093 -83 1127
rect -117 1025 -83 1059
rect -117 957 -83 991
rect -117 889 -83 923
rect -117 821 -83 855
rect -117 753 -83 787
rect -117 685 -83 719
rect -117 617 -83 651
rect -117 549 -83 583
rect -117 481 -83 515
rect -117 413 -83 447
rect -117 345 -83 379
rect -117 277 -83 311
rect -117 209 -83 243
rect -117 141 -83 175
rect -117 73 -83 107
rect -117 5 -83 39
rect -117 -63 -83 -29
rect -117 -131 -83 -97
rect -117 -199 -83 -165
rect -117 -267 -83 -233
rect -117 -343 -83 -301
rect 3993 9661 4027 9703
rect 3993 9593 4027 9627
rect 3993 9525 4027 9559
rect 3993 9457 4027 9491
rect 3993 9389 4027 9423
rect 3993 9321 4027 9355
rect 3993 9253 4027 9287
rect 3993 9185 4027 9219
rect 3993 9117 4027 9151
rect 3993 9049 4027 9083
rect 3993 8981 4027 9015
rect 3993 8913 4027 8947
rect 3993 8845 4027 8879
rect 3993 8777 4027 8811
rect 3993 8709 4027 8743
rect 3993 8641 4027 8675
rect 3993 8573 4027 8607
rect 3993 8505 4027 8539
rect 3993 8437 4027 8471
rect 3993 8369 4027 8403
rect 3993 8301 4027 8335
rect 3993 8233 4027 8267
rect 3993 8165 4027 8199
rect 3993 8097 4027 8131
rect 3993 8029 4027 8063
rect 3993 7961 4027 7995
rect 3993 7893 4027 7927
rect 3993 7825 4027 7859
rect 3993 7757 4027 7791
rect 3993 7689 4027 7723
rect 3993 7621 4027 7655
rect 3993 7553 4027 7587
rect 3993 7485 4027 7519
rect 3993 7417 4027 7451
rect 3993 7349 4027 7383
rect 3993 7281 4027 7315
rect 3993 7213 4027 7247
rect 3993 7145 4027 7179
rect 3993 7077 4027 7111
rect 3993 7009 4027 7043
rect 3993 6941 4027 6975
rect 3993 6873 4027 6907
rect 3993 6805 4027 6839
rect 3993 6737 4027 6771
rect 3993 6669 4027 6703
rect 3993 6601 4027 6635
rect 3993 6533 4027 6567
rect 3993 6465 4027 6499
rect 3993 6397 4027 6431
rect 3993 6329 4027 6363
rect 3993 6261 4027 6295
rect 3993 6193 4027 6227
rect 3993 6125 4027 6159
rect 3993 6057 4027 6091
rect 3993 5989 4027 6023
rect 3993 5921 4027 5955
rect 3993 5853 4027 5887
rect 3993 5785 4027 5819
rect 3993 5717 4027 5751
rect 3993 5649 4027 5683
rect 3993 5581 4027 5615
rect 3993 5513 4027 5547
rect 3993 5445 4027 5479
rect 3993 5377 4027 5411
rect 3993 5309 4027 5343
rect 3993 5241 4027 5275
rect 3993 5173 4027 5207
rect 3993 5105 4027 5139
rect 3993 5037 4027 5071
rect 3993 4969 4027 5003
rect 3993 4901 4027 4935
rect 3993 4833 4027 4867
rect 3993 4765 4027 4799
rect 3993 4697 4027 4731
rect 3993 4629 4027 4663
rect 3993 4561 4027 4595
rect 3993 4493 4027 4527
rect 3993 4425 4027 4459
rect 3993 4357 4027 4391
rect 3993 4289 4027 4323
rect 3993 4221 4027 4255
rect 3993 4153 4027 4187
rect 3993 4085 4027 4119
rect 3993 4017 4027 4051
rect 3993 3949 4027 3983
rect 3993 3881 4027 3915
rect 3993 3813 4027 3847
rect 3993 3745 4027 3779
rect 3993 3677 4027 3711
rect 3993 3609 4027 3643
rect 3993 3541 4027 3575
rect 3993 3473 4027 3507
rect 3993 3405 4027 3439
rect 3993 3337 4027 3371
rect 3993 3269 4027 3303
rect 3993 3201 4027 3235
rect 3993 3133 4027 3167
rect 3993 3065 4027 3099
rect 3993 2997 4027 3031
rect 3993 2929 4027 2963
rect 3993 2861 4027 2895
rect 3993 2793 4027 2827
rect 3993 2725 4027 2759
rect 3993 2657 4027 2691
rect 3993 2589 4027 2623
rect 3993 2521 4027 2555
rect 3993 2453 4027 2487
rect 3993 2385 4027 2419
rect 3993 2317 4027 2351
rect 3993 2249 4027 2283
rect 3993 2181 4027 2215
rect 3993 2113 4027 2147
rect 3993 2045 4027 2079
rect 3993 1977 4027 2011
rect 3993 1909 4027 1943
rect 3993 1841 4027 1875
rect 3993 1773 4027 1807
rect 3993 1705 4027 1739
rect 3993 1637 4027 1671
rect 3993 1569 4027 1603
rect 3993 1501 4027 1535
rect 3993 1433 4027 1467
rect 3993 1365 4027 1399
rect 3993 1297 4027 1331
rect 3993 1229 4027 1263
rect 3993 1161 4027 1195
rect 3993 1093 4027 1127
rect 3993 1025 4027 1059
rect 3993 957 4027 991
rect 3993 889 4027 923
rect 3993 821 4027 855
rect 3993 753 4027 787
rect 3993 685 4027 719
rect 3993 617 4027 651
rect 3993 549 4027 583
rect 3993 481 4027 515
rect 3993 413 4027 447
rect 3993 345 4027 379
rect 3993 277 4027 311
rect 3993 209 4027 243
rect 3993 141 4027 175
rect 3993 73 4027 107
rect 3993 5 4027 39
rect 3993 -63 4027 -29
rect 3993 -131 4027 -97
rect 3993 -199 4027 -165
rect 3993 -267 4027 -233
rect 3993 -343 4027 -301
rect -117 -377 -34 -343
rect 0 -377 34 -343
rect 68 -377 102 -343
rect 136 -377 170 -343
rect 204 -377 238 -343
rect 272 -377 306 -343
rect 340 -377 374 -343
rect 408 -377 442 -343
rect 476 -377 510 -343
rect 544 -377 578 -343
rect 612 -377 646 -343
rect 680 -377 714 -343
rect 748 -377 782 -343
rect 816 -377 850 -343
rect 884 -377 918 -343
rect 952 -377 986 -343
rect 1020 -377 1054 -343
rect 1088 -377 1122 -343
rect 1156 -377 1190 -343
rect 1224 -377 1258 -343
rect 1292 -377 1326 -343
rect 1360 -377 1394 -343
rect 1428 -377 1462 -343
rect 1496 -377 1530 -343
rect 1564 -377 1598 -343
rect 1632 -377 1666 -343
rect 1700 -377 1734 -343
rect 1768 -377 1802 -343
rect 1836 -377 1870 -343
rect 1904 -377 1938 -343
rect 1972 -377 2006 -343
rect 2040 -377 2074 -343
rect 2108 -377 2142 -343
rect 2176 -377 2210 -343
rect 2244 -377 2278 -343
rect 2312 -377 2346 -343
rect 2380 -377 2414 -343
rect 2448 -377 2482 -343
rect 2516 -377 2550 -343
rect 2584 -377 2618 -343
rect 2652 -377 2686 -343
rect 2720 -377 2754 -343
rect 2788 -377 2822 -343
rect 2856 -377 2890 -343
rect 2924 -377 2958 -343
rect 2992 -377 3026 -343
rect 3060 -377 3094 -343
rect 3128 -377 3162 -343
rect 3196 -377 3230 -343
rect 3264 -377 3298 -343
rect 3332 -377 3366 -343
rect 3400 -377 3434 -343
rect 3468 -377 3502 -343
rect 3536 -377 3570 -343
rect 3604 -377 3638 -343
rect 3672 -377 3706 -343
rect 3740 -377 3774 -343
rect 3808 -377 3842 -343
rect 3876 -377 3910 -343
rect 3944 -377 4027 -343
<< metal1 >>
rect 170 9420 3790 9630
rect 170 9356 460 9420
rect 170 9304 204 9356
rect 256 9304 284 9356
rect 336 9304 460 9356
rect 170 8186 460 9304
rect 560 9356 720 9360
rect 560 9304 574 9356
rect 626 9304 654 9356
rect 706 9304 720 9356
rect 560 9300 720 9304
rect 930 9356 1090 9360
rect 930 9304 944 9356
rect 996 9304 1024 9356
rect 1076 9304 1090 9356
rect 930 9300 1090 9304
rect 1300 9356 1460 9360
rect 1300 9304 1314 9356
rect 1366 9304 1394 9356
rect 1446 9304 1460 9356
rect 1300 9300 1460 9304
rect 1670 9356 1830 9360
rect 1670 9304 1684 9356
rect 1736 9304 1764 9356
rect 1816 9304 1830 9356
rect 1670 9300 1830 9304
rect 2040 9356 2200 9360
rect 2040 9304 2054 9356
rect 2106 9304 2134 9356
rect 2186 9304 2200 9356
rect 2040 9300 2200 9304
rect 2410 9356 2570 9360
rect 2410 9304 2424 9356
rect 2476 9304 2504 9356
rect 2556 9304 2570 9356
rect 2410 9300 2570 9304
rect 2780 9356 2940 9360
rect 2780 9304 2794 9356
rect 2846 9304 2874 9356
rect 2926 9304 2940 9356
rect 2780 9300 2940 9304
rect 3150 9356 3310 9360
rect 3150 9304 3164 9356
rect 3216 9304 3244 9356
rect 3296 9304 3310 9356
rect 3150 9300 3310 9304
rect 3500 9356 3790 9420
rect 3500 9304 3534 9356
rect 3586 9304 3614 9356
rect 3666 9304 3790 9356
rect 770 8310 830 9160
rect 1140 8310 1200 9160
rect 1510 8310 1570 9160
rect 1880 8310 1940 9160
rect 2250 8310 2310 9160
rect 2620 8310 2680 9160
rect 2990 8310 3050 9160
rect 3360 8310 3420 9160
rect 540 8306 830 8310
rect 540 8254 574 8306
rect 626 8254 654 8306
rect 706 8254 830 8306
rect 540 8250 830 8254
rect 910 8306 1200 8310
rect 910 8254 944 8306
rect 996 8254 1024 8306
rect 1076 8254 1200 8306
rect 910 8250 1200 8254
rect 1280 8306 1570 8310
rect 1280 8254 1314 8306
rect 1366 8254 1394 8306
rect 1446 8254 1570 8306
rect 1280 8250 1570 8254
rect 1650 8306 1940 8310
rect 1650 8254 1684 8306
rect 1736 8254 1764 8306
rect 1816 8254 1940 8306
rect 1650 8250 1940 8254
rect 2020 8306 2310 8310
rect 2020 8254 2054 8306
rect 2106 8254 2134 8306
rect 2186 8254 2310 8306
rect 2020 8250 2310 8254
rect 2390 8306 2680 8310
rect 2390 8254 2424 8306
rect 2476 8254 2504 8306
rect 2556 8254 2680 8306
rect 2390 8250 2680 8254
rect 2760 8306 3050 8310
rect 2760 8254 2794 8306
rect 2846 8254 2874 8306
rect 2926 8254 3050 8306
rect 2760 8250 3050 8254
rect 3130 8306 3420 8310
rect 3130 8254 3164 8306
rect 3216 8254 3244 8306
rect 3296 8254 3420 8306
rect 3130 8250 3420 8254
rect 170 8134 204 8186
rect 256 8134 284 8186
rect 336 8134 460 8186
rect 170 7016 460 8134
rect 560 8186 720 8190
rect 560 8134 574 8186
rect 626 8134 654 8186
rect 706 8134 720 8186
rect 560 8130 720 8134
rect 930 8186 1090 8190
rect 930 8134 944 8186
rect 996 8134 1024 8186
rect 1076 8134 1090 8186
rect 930 8130 1090 8134
rect 1300 8186 1460 8190
rect 1300 8134 1314 8186
rect 1366 8134 1394 8186
rect 1446 8134 1460 8186
rect 1300 8130 1460 8134
rect 1670 8186 1830 8190
rect 1670 8134 1684 8186
rect 1736 8134 1764 8186
rect 1816 8134 1830 8186
rect 1670 8130 1830 8134
rect 2040 8186 2200 8190
rect 2040 8134 2054 8186
rect 2106 8134 2134 8186
rect 2186 8134 2200 8186
rect 2040 8130 2200 8134
rect 2410 8186 2570 8190
rect 2410 8134 2424 8186
rect 2476 8134 2504 8186
rect 2556 8134 2570 8186
rect 2410 8130 2570 8134
rect 2780 8186 2940 8190
rect 2780 8134 2794 8186
rect 2846 8134 2874 8186
rect 2926 8134 2940 8186
rect 2780 8130 2940 8134
rect 3150 8186 3310 8190
rect 3150 8134 3164 8186
rect 3216 8134 3244 8186
rect 3296 8134 3310 8186
rect 3150 8130 3310 8134
rect 3500 8186 3790 9304
rect 3500 8134 3534 8186
rect 3586 8134 3614 8186
rect 3666 8134 3790 8186
rect 770 7140 830 7990
rect 1140 7140 1200 7990
rect 1510 7140 1570 7990
rect 1880 7140 1940 7990
rect 2250 7140 2310 7990
rect 2620 7140 2680 7990
rect 2990 7140 3050 7990
rect 3360 7140 3420 7990
rect 540 7136 830 7140
rect 540 7084 574 7136
rect 626 7084 654 7136
rect 706 7084 830 7136
rect 540 7080 830 7084
rect 910 7136 1200 7140
rect 910 7084 944 7136
rect 996 7084 1024 7136
rect 1076 7084 1200 7136
rect 910 7080 1200 7084
rect 1280 7136 1570 7140
rect 1280 7084 1314 7136
rect 1366 7084 1394 7136
rect 1446 7084 1570 7136
rect 1280 7080 1570 7084
rect 1650 7136 1940 7140
rect 1650 7084 1684 7136
rect 1736 7084 1764 7136
rect 1816 7084 1940 7136
rect 1650 7080 1940 7084
rect 2020 7136 2310 7140
rect 2020 7084 2054 7136
rect 2106 7084 2134 7136
rect 2186 7084 2310 7136
rect 2020 7080 2310 7084
rect 2390 7136 2680 7140
rect 2390 7084 2424 7136
rect 2476 7084 2504 7136
rect 2556 7084 2680 7136
rect 2390 7080 2680 7084
rect 2760 7136 3050 7140
rect 2760 7084 2794 7136
rect 2846 7084 2874 7136
rect 2926 7084 3050 7136
rect 2760 7080 3050 7084
rect 3130 7136 3420 7140
rect 3130 7084 3164 7136
rect 3216 7084 3244 7136
rect 3296 7084 3420 7136
rect 3130 7080 3420 7084
rect 170 6964 204 7016
rect 256 6964 284 7016
rect 336 6964 460 7016
rect 170 5846 460 6964
rect 560 7016 720 7020
rect 560 6964 574 7016
rect 626 6964 654 7016
rect 706 6964 720 7016
rect 560 6960 720 6964
rect 930 7016 1090 7020
rect 930 6964 944 7016
rect 996 6964 1024 7016
rect 1076 6964 1090 7016
rect 930 6960 1090 6964
rect 1300 7016 1460 7020
rect 1300 6964 1314 7016
rect 1366 6964 1394 7016
rect 1446 6964 1460 7016
rect 1300 6960 1460 6964
rect 1670 7016 1830 7020
rect 1670 6964 1684 7016
rect 1736 6964 1764 7016
rect 1816 6964 1830 7016
rect 1670 6960 1830 6964
rect 2040 7016 2200 7020
rect 2040 6964 2054 7016
rect 2106 6964 2134 7016
rect 2186 6964 2200 7016
rect 2040 6960 2200 6964
rect 2410 7016 2570 7020
rect 2410 6964 2424 7016
rect 2476 6964 2504 7016
rect 2556 6964 2570 7016
rect 2410 6960 2570 6964
rect 2780 7016 2940 7020
rect 2780 6964 2794 7016
rect 2846 6964 2874 7016
rect 2926 6964 2940 7016
rect 2780 6960 2940 6964
rect 3150 7016 3310 7020
rect 3150 6964 3164 7016
rect 3216 6964 3244 7016
rect 3296 6964 3310 7016
rect 3150 6960 3310 6964
rect 3500 7016 3790 8134
rect 3500 6964 3534 7016
rect 3586 6964 3614 7016
rect 3666 6964 3790 7016
rect 770 5970 830 6820
rect 1140 5970 1200 6820
rect 1510 5970 1570 6820
rect 1880 5970 1940 6820
rect 2250 5970 2310 6820
rect 2620 5970 2680 6820
rect 2990 5970 3050 6820
rect 3360 5970 3420 6820
rect 540 5966 830 5970
rect 540 5914 574 5966
rect 626 5914 654 5966
rect 706 5914 830 5966
rect 540 5910 830 5914
rect 910 5966 1200 5970
rect 910 5914 944 5966
rect 996 5914 1024 5966
rect 1076 5914 1200 5966
rect 910 5910 1200 5914
rect 1280 5966 1570 5970
rect 1280 5914 1314 5966
rect 1366 5914 1394 5966
rect 1446 5914 1570 5966
rect 1280 5910 1570 5914
rect 1650 5966 1940 5970
rect 1650 5914 1684 5966
rect 1736 5914 1764 5966
rect 1816 5914 1940 5966
rect 1650 5910 1940 5914
rect 2020 5966 2310 5970
rect 2020 5914 2054 5966
rect 2106 5914 2134 5966
rect 2186 5914 2310 5966
rect 2020 5910 2310 5914
rect 2390 5966 2680 5970
rect 2390 5914 2424 5966
rect 2476 5914 2504 5966
rect 2556 5914 2680 5966
rect 2390 5910 2680 5914
rect 2760 5966 3050 5970
rect 2760 5914 2794 5966
rect 2846 5914 2874 5966
rect 2926 5914 3050 5966
rect 2760 5910 3050 5914
rect 3130 5966 3420 5970
rect 3130 5914 3164 5966
rect 3216 5914 3244 5966
rect 3296 5914 3420 5966
rect 3130 5910 3420 5914
rect 170 5794 204 5846
rect 256 5794 284 5846
rect 336 5794 460 5846
rect 170 4616 460 5794
rect 560 5846 720 5850
rect 560 5794 574 5846
rect 626 5794 654 5846
rect 706 5794 720 5846
rect 560 5790 720 5794
rect 930 5846 1090 5850
rect 930 5794 944 5846
rect 996 5794 1024 5846
rect 1076 5794 1090 5846
rect 930 5790 1090 5794
rect 1300 5846 1460 5850
rect 1300 5794 1314 5846
rect 1366 5794 1394 5846
rect 1446 5794 1460 5846
rect 1300 5790 1460 5794
rect 1670 5846 1830 5850
rect 1670 5794 1684 5846
rect 1736 5794 1764 5846
rect 1816 5794 1830 5846
rect 1670 5790 1830 5794
rect 2040 5846 2320 5850
rect 2040 5794 2054 5846
rect 2106 5794 2134 5846
rect 2186 5794 2320 5846
rect 2040 5790 2320 5794
rect 2410 5846 2570 5850
rect 2410 5794 2424 5846
rect 2476 5794 2504 5846
rect 2556 5794 2570 5846
rect 2410 5790 2570 5794
rect 2780 5846 2940 5850
rect 2780 5794 2794 5846
rect 2846 5794 2874 5846
rect 2926 5794 2940 5846
rect 2780 5790 2940 5794
rect 3150 5846 3310 5850
rect 3150 5794 3164 5846
rect 3216 5794 3244 5846
rect 3296 5794 3310 5846
rect 3150 5790 3310 5794
rect 3500 5846 3790 6964
rect 3500 5794 3534 5846
rect 3586 5794 3614 5846
rect 3666 5794 3790 5846
rect 2250 5650 2320 5790
rect 770 4800 830 5650
rect 1140 4800 1200 5650
rect 1510 4800 1570 5650
rect 1880 5101 1940 5650
rect 1880 5049 1884 5101
rect 1936 5049 1940 5101
rect 1880 5011 1940 5049
rect 1880 4959 1884 5011
rect 1936 4959 1940 5011
rect 1880 4940 1940 4959
rect 2250 4800 2310 5650
rect 2620 4800 2680 5650
rect 2990 4800 3050 5650
rect 3360 4800 3420 5650
rect 540 4796 830 4800
rect 540 4744 574 4796
rect 626 4744 654 4796
rect 706 4744 830 4796
rect 540 4740 830 4744
rect 910 4796 1200 4800
rect 910 4744 944 4796
rect 996 4744 1024 4796
rect 1076 4744 1200 4796
rect 910 4740 1200 4744
rect 1280 4796 1570 4800
rect 1280 4744 1314 4796
rect 1366 4744 1394 4796
rect 1446 4744 1570 4796
rect 1280 4740 1570 4744
rect 1670 4710 1830 4800
rect 2050 4740 2310 4800
rect 2390 4796 2680 4800
rect 2390 4744 2424 4796
rect 2476 4744 2504 4796
rect 2556 4744 2680 4796
rect 2390 4740 2680 4744
rect 2760 4796 3050 4800
rect 2760 4744 2794 4796
rect 2846 4744 2874 4796
rect 2926 4744 3050 4796
rect 2760 4740 3050 4744
rect 3130 4796 3420 4800
rect 3130 4744 3164 4796
rect 3216 4744 3244 4796
rect 3296 4744 3420 4796
rect 3130 4740 3420 4744
rect 1670 4706 2020 4710
rect 1670 4654 1704 4706
rect 1756 4654 1804 4706
rect 1856 4654 1904 4706
rect 1956 4654 2020 4706
rect 1670 4650 2020 4654
rect 170 4564 204 4616
rect 256 4564 284 4616
rect 336 4564 460 4616
rect 170 3446 460 4564
rect 560 4616 720 4620
rect 560 4564 574 4616
rect 626 4564 654 4616
rect 706 4564 720 4616
rect 560 4560 720 4564
rect 930 4616 1090 4620
rect 930 4564 944 4616
rect 996 4564 1024 4616
rect 1076 4564 1090 4616
rect 930 4560 1090 4564
rect 1300 4616 1460 4620
rect 1300 4564 1314 4616
rect 1366 4564 1394 4616
rect 1446 4564 1460 4616
rect 1300 4560 1460 4564
rect 1670 4616 1940 4620
rect 1670 4564 1684 4616
rect 1736 4564 1764 4616
rect 1816 4564 1940 4616
rect 1670 4560 1940 4564
rect 770 3570 830 4420
rect 1140 3570 1200 4420
rect 1510 3570 1570 4420
rect 1880 3570 1940 4560
rect 540 3566 830 3570
rect 540 3514 574 3566
rect 626 3514 654 3566
rect 706 3514 830 3566
rect 540 3510 830 3514
rect 910 3566 1200 3570
rect 910 3514 944 3566
rect 996 3514 1024 3566
rect 1076 3514 1200 3566
rect 910 3510 1200 3514
rect 1280 3566 1570 3570
rect 1280 3514 1314 3566
rect 1366 3514 1394 3566
rect 1446 3514 1570 3566
rect 1280 3510 1570 3514
rect 1650 3510 1940 3570
rect 1970 3570 2020 4650
rect 2120 4616 2200 4620
rect 2120 4564 2134 4616
rect 2186 4564 2200 4616
rect 2120 4560 2200 4564
rect 2410 4616 2570 4620
rect 2410 4564 2424 4616
rect 2476 4564 2504 4616
rect 2556 4564 2570 4616
rect 2410 4560 2570 4564
rect 2780 4616 2940 4620
rect 2780 4564 2794 4616
rect 2846 4564 2874 4616
rect 2926 4564 2940 4616
rect 2780 4560 2940 4564
rect 3150 4616 3310 4620
rect 3150 4564 3164 4616
rect 3216 4564 3244 4616
rect 3296 4564 3310 4616
rect 3150 4560 3310 4564
rect 3500 4616 3790 5794
rect 3500 4564 3534 4616
rect 3586 4564 3614 4616
rect 3666 4564 3790 4616
rect 2250 3856 2310 4420
rect 2250 3804 2254 3856
rect 2306 3804 2310 3856
rect 2250 3776 2310 3804
rect 2250 3724 2254 3776
rect 2306 3724 2310 3776
rect 2250 3710 2310 3724
rect 2620 3570 2680 4420
rect 2990 3570 3050 4420
rect 3360 3570 3420 4420
rect 1970 3510 2200 3570
rect 2390 3566 2680 3570
rect 2390 3514 2424 3566
rect 2476 3514 2504 3566
rect 2556 3514 2680 3566
rect 2390 3510 2680 3514
rect 2760 3566 3050 3570
rect 2760 3514 2794 3566
rect 2846 3514 2874 3566
rect 2926 3514 3050 3566
rect 2760 3510 3050 3514
rect 3130 3566 3420 3570
rect 3130 3514 3164 3566
rect 3216 3514 3244 3566
rect 3296 3514 3420 3566
rect 3130 3510 3420 3514
rect 170 3394 204 3446
rect 256 3394 284 3446
rect 336 3394 460 3446
rect 170 2276 460 3394
rect 560 3446 720 3450
rect 560 3394 574 3446
rect 626 3394 654 3446
rect 706 3394 720 3446
rect 560 3390 720 3394
rect 930 3446 1090 3450
rect 930 3394 944 3446
rect 996 3394 1024 3446
rect 1076 3394 1090 3446
rect 930 3390 1090 3394
rect 1300 3446 1460 3450
rect 1300 3394 1314 3446
rect 1366 3394 1394 3446
rect 1446 3394 1460 3446
rect 1300 3390 1460 3394
rect 1670 3446 1830 3450
rect 1670 3394 1684 3446
rect 1736 3394 1764 3446
rect 1816 3394 1830 3446
rect 1670 3390 1830 3394
rect 2040 3446 2200 3450
rect 2040 3394 2054 3446
rect 2106 3394 2134 3446
rect 2186 3394 2200 3446
rect 2040 3390 2200 3394
rect 2410 3446 2570 3450
rect 2410 3394 2424 3446
rect 2476 3394 2504 3446
rect 2556 3394 2570 3446
rect 2410 3390 2570 3394
rect 2780 3446 2940 3450
rect 2780 3394 2794 3446
rect 2846 3394 2874 3446
rect 2926 3394 2940 3446
rect 2780 3390 2940 3394
rect 3150 3446 3310 3450
rect 3150 3394 3164 3446
rect 3216 3394 3244 3446
rect 3296 3394 3310 3446
rect 3150 3390 3310 3394
rect 3500 3446 3790 4564
rect 3500 3394 3534 3446
rect 3586 3394 3614 3446
rect 3666 3394 3790 3446
rect 770 2400 830 3250
rect 1140 2400 1200 3250
rect 1510 2400 1570 3250
rect 1880 2400 1940 3250
rect 2250 2400 2310 3250
rect 2620 2400 2680 3250
rect 2990 2400 3050 3250
rect 3360 2400 3420 3250
rect 540 2396 830 2400
rect 540 2344 574 2396
rect 626 2344 654 2396
rect 706 2344 830 2396
rect 540 2340 830 2344
rect 910 2396 1200 2400
rect 910 2344 944 2396
rect 996 2344 1024 2396
rect 1076 2344 1200 2396
rect 910 2340 1200 2344
rect 1280 2396 1570 2400
rect 1280 2344 1314 2396
rect 1366 2344 1394 2396
rect 1446 2344 1570 2396
rect 1280 2340 1570 2344
rect 1650 2396 1940 2400
rect 1650 2344 1684 2396
rect 1736 2344 1764 2396
rect 1816 2344 1940 2396
rect 1650 2340 1940 2344
rect 2020 2396 2310 2400
rect 2020 2344 2054 2396
rect 2106 2344 2134 2396
rect 2186 2344 2310 2396
rect 2020 2340 2310 2344
rect 2390 2396 2680 2400
rect 2390 2344 2424 2396
rect 2476 2344 2504 2396
rect 2556 2344 2680 2396
rect 2390 2340 2680 2344
rect 2760 2396 3050 2400
rect 2760 2344 2794 2396
rect 2846 2344 2874 2396
rect 2926 2344 3050 2396
rect 2760 2340 3050 2344
rect 3130 2396 3420 2400
rect 3130 2344 3164 2396
rect 3216 2344 3244 2396
rect 3296 2344 3420 2396
rect 3130 2340 3420 2344
rect 170 2224 204 2276
rect 256 2224 284 2276
rect 336 2224 460 2276
rect 170 1106 460 2224
rect 560 2276 720 2280
rect 560 2224 574 2276
rect 626 2224 654 2276
rect 706 2224 720 2276
rect 560 2220 720 2224
rect 930 2276 1090 2280
rect 930 2224 944 2276
rect 996 2224 1024 2276
rect 1076 2224 1090 2276
rect 930 2220 1090 2224
rect 1300 2276 1460 2280
rect 1300 2224 1314 2276
rect 1366 2224 1394 2276
rect 1446 2224 1460 2276
rect 1300 2220 1460 2224
rect 1670 2276 1830 2280
rect 1670 2224 1684 2276
rect 1736 2224 1764 2276
rect 1816 2224 1830 2276
rect 1670 2220 1830 2224
rect 2040 2276 2200 2280
rect 2040 2224 2054 2276
rect 2106 2224 2134 2276
rect 2186 2224 2200 2276
rect 2040 2220 2200 2224
rect 2410 2276 2570 2280
rect 2410 2224 2424 2276
rect 2476 2224 2504 2276
rect 2556 2224 2570 2276
rect 2410 2220 2570 2224
rect 2780 2276 2940 2280
rect 2780 2224 2794 2276
rect 2846 2224 2874 2276
rect 2926 2224 2940 2276
rect 2780 2220 2940 2224
rect 3150 2276 3310 2280
rect 3150 2224 3164 2276
rect 3216 2224 3244 2276
rect 3296 2224 3310 2276
rect 3150 2220 3310 2224
rect 3500 2276 3790 3394
rect 3500 2224 3534 2276
rect 3586 2224 3614 2276
rect 3666 2224 3790 2276
rect 770 1230 830 2080
rect 1140 1230 1200 2080
rect 1510 1230 1570 2080
rect 1880 1230 1940 2080
rect 2250 1230 2310 2080
rect 2620 1230 2680 2080
rect 2990 1230 3050 2080
rect 3360 1230 3420 2080
rect 540 1226 830 1230
rect 540 1174 574 1226
rect 626 1174 654 1226
rect 706 1174 830 1226
rect 540 1170 830 1174
rect 910 1226 1200 1230
rect 910 1174 944 1226
rect 996 1174 1024 1226
rect 1076 1174 1200 1226
rect 910 1170 1200 1174
rect 1280 1226 1570 1230
rect 1280 1174 1314 1226
rect 1366 1174 1394 1226
rect 1446 1174 1570 1226
rect 1280 1170 1570 1174
rect 1650 1226 1940 1230
rect 1650 1174 1684 1226
rect 1736 1174 1764 1226
rect 1816 1174 1940 1226
rect 1650 1170 1940 1174
rect 2020 1226 2310 1230
rect 2020 1174 2054 1226
rect 2106 1174 2134 1226
rect 2186 1174 2310 1226
rect 2020 1170 2310 1174
rect 2390 1226 2680 1230
rect 2390 1174 2424 1226
rect 2476 1174 2504 1226
rect 2556 1174 2680 1226
rect 2390 1170 2680 1174
rect 2760 1226 3050 1230
rect 2760 1174 2794 1226
rect 2846 1174 2874 1226
rect 2926 1174 3050 1226
rect 2760 1170 3050 1174
rect 3130 1226 3420 1230
rect 3130 1174 3164 1226
rect 3216 1174 3244 1226
rect 3296 1174 3420 1226
rect 3130 1170 3420 1174
rect 170 1054 204 1106
rect 256 1054 284 1106
rect 336 1054 460 1106
rect 170 -60 460 1054
rect 560 1106 720 1110
rect 560 1054 574 1106
rect 626 1054 654 1106
rect 706 1054 720 1106
rect 560 1050 720 1054
rect 930 1106 1090 1110
rect 930 1054 944 1106
rect 996 1054 1024 1106
rect 1076 1054 1090 1106
rect 930 1050 1090 1054
rect 1300 1106 1460 1110
rect 1300 1054 1314 1106
rect 1366 1054 1394 1106
rect 1446 1054 1460 1106
rect 1300 1050 1460 1054
rect 1670 1106 1830 1110
rect 1670 1054 1684 1106
rect 1736 1054 1764 1106
rect 1816 1054 1830 1106
rect 1670 1050 1830 1054
rect 2040 1106 2200 1110
rect 2040 1054 2054 1106
rect 2106 1054 2134 1106
rect 2186 1054 2200 1106
rect 2040 1050 2200 1054
rect 2410 1106 2570 1110
rect 2410 1054 2424 1106
rect 2476 1054 2504 1106
rect 2556 1054 2570 1106
rect 2410 1050 2570 1054
rect 2780 1106 2940 1110
rect 2780 1054 2794 1106
rect 2846 1054 2874 1106
rect 2926 1054 2940 1106
rect 2780 1050 2940 1054
rect 3150 1106 3310 1110
rect 3150 1054 3164 1106
rect 3216 1054 3244 1106
rect 3296 1054 3310 1106
rect 3150 1050 3310 1054
rect 3500 1106 3790 2224
rect 3500 1054 3534 1106
rect 3586 1054 3614 1106
rect 3666 1054 3790 1106
rect 770 60 830 910
rect 1140 60 1200 910
rect 1510 60 1570 910
rect 1880 60 1940 910
rect 2250 60 2310 910
rect 2620 60 2680 910
rect 2990 60 3050 910
rect 3360 60 3420 910
rect 540 56 830 60
rect 540 4 574 56
rect 626 4 654 56
rect 706 4 830 56
rect 540 0 830 4
rect 910 56 1200 60
rect 910 4 944 56
rect 996 4 1024 56
rect 1076 4 1200 56
rect 910 0 1200 4
rect 1280 56 1570 60
rect 1280 4 1314 56
rect 1366 4 1394 56
rect 1446 4 1570 56
rect 1280 0 1570 4
rect 1650 56 1940 60
rect 1650 4 1684 56
rect 1736 4 1764 56
rect 1816 4 1940 56
rect 1650 0 1940 4
rect 2020 56 2310 60
rect 2020 4 2054 56
rect 2106 4 2134 56
rect 2186 4 2310 56
rect 2020 0 2310 4
rect 2390 56 2680 60
rect 2390 4 2424 56
rect 2476 4 2504 56
rect 2556 4 2680 56
rect 2390 0 2680 4
rect 2760 56 3050 60
rect 2760 4 2794 56
rect 2846 4 2874 56
rect 2926 4 3050 56
rect 2760 0 3050 4
rect 3130 56 3420 60
rect 3130 4 3164 56
rect 3216 4 3244 56
rect 3296 4 3420 56
rect 3130 0 3420 4
rect 3500 -60 3790 1054
rect 170 -270 3790 -60
<< via1 >>
rect 204 9304 256 9356
rect 284 9304 336 9356
rect 574 9304 626 9356
rect 654 9304 706 9356
rect 944 9304 996 9356
rect 1024 9304 1076 9356
rect 1314 9304 1366 9356
rect 1394 9304 1446 9356
rect 1684 9304 1736 9356
rect 1764 9304 1816 9356
rect 2054 9304 2106 9356
rect 2134 9304 2186 9356
rect 2424 9304 2476 9356
rect 2504 9304 2556 9356
rect 2794 9304 2846 9356
rect 2874 9304 2926 9356
rect 3164 9304 3216 9356
rect 3244 9304 3296 9356
rect 3534 9304 3586 9356
rect 3614 9304 3666 9356
rect 574 8254 626 8306
rect 654 8254 706 8306
rect 944 8254 996 8306
rect 1024 8254 1076 8306
rect 1314 8254 1366 8306
rect 1394 8254 1446 8306
rect 1684 8254 1736 8306
rect 1764 8254 1816 8306
rect 2054 8254 2106 8306
rect 2134 8254 2186 8306
rect 2424 8254 2476 8306
rect 2504 8254 2556 8306
rect 2794 8254 2846 8306
rect 2874 8254 2926 8306
rect 3164 8254 3216 8306
rect 3244 8254 3296 8306
rect 204 8134 256 8186
rect 284 8134 336 8186
rect 574 8134 626 8186
rect 654 8134 706 8186
rect 944 8134 996 8186
rect 1024 8134 1076 8186
rect 1314 8134 1366 8186
rect 1394 8134 1446 8186
rect 1684 8134 1736 8186
rect 1764 8134 1816 8186
rect 2054 8134 2106 8186
rect 2134 8134 2186 8186
rect 2424 8134 2476 8186
rect 2504 8134 2556 8186
rect 2794 8134 2846 8186
rect 2874 8134 2926 8186
rect 3164 8134 3216 8186
rect 3244 8134 3296 8186
rect 3534 8134 3586 8186
rect 3614 8134 3666 8186
rect 574 7084 626 7136
rect 654 7084 706 7136
rect 944 7084 996 7136
rect 1024 7084 1076 7136
rect 1314 7084 1366 7136
rect 1394 7084 1446 7136
rect 1684 7084 1736 7136
rect 1764 7084 1816 7136
rect 2054 7084 2106 7136
rect 2134 7084 2186 7136
rect 2424 7084 2476 7136
rect 2504 7084 2556 7136
rect 2794 7084 2846 7136
rect 2874 7084 2926 7136
rect 3164 7084 3216 7136
rect 3244 7084 3296 7136
rect 204 6964 256 7016
rect 284 6964 336 7016
rect 574 6964 626 7016
rect 654 6964 706 7016
rect 944 6964 996 7016
rect 1024 6964 1076 7016
rect 1314 6964 1366 7016
rect 1394 6964 1446 7016
rect 1684 6964 1736 7016
rect 1764 6964 1816 7016
rect 2054 6964 2106 7016
rect 2134 6964 2186 7016
rect 2424 6964 2476 7016
rect 2504 6964 2556 7016
rect 2794 6964 2846 7016
rect 2874 6964 2926 7016
rect 3164 6964 3216 7016
rect 3244 6964 3296 7016
rect 3534 6964 3586 7016
rect 3614 6964 3666 7016
rect 574 5914 626 5966
rect 654 5914 706 5966
rect 944 5914 996 5966
rect 1024 5914 1076 5966
rect 1314 5914 1366 5966
rect 1394 5914 1446 5966
rect 1684 5914 1736 5966
rect 1764 5914 1816 5966
rect 2054 5914 2106 5966
rect 2134 5914 2186 5966
rect 2424 5914 2476 5966
rect 2504 5914 2556 5966
rect 2794 5914 2846 5966
rect 2874 5914 2926 5966
rect 3164 5914 3216 5966
rect 3244 5914 3296 5966
rect 204 5794 256 5846
rect 284 5794 336 5846
rect 574 5794 626 5846
rect 654 5794 706 5846
rect 944 5794 996 5846
rect 1024 5794 1076 5846
rect 1314 5794 1366 5846
rect 1394 5794 1446 5846
rect 1684 5794 1736 5846
rect 1764 5794 1816 5846
rect 2054 5794 2106 5846
rect 2134 5794 2186 5846
rect 2424 5794 2476 5846
rect 2504 5794 2556 5846
rect 2794 5794 2846 5846
rect 2874 5794 2926 5846
rect 3164 5794 3216 5846
rect 3244 5794 3296 5846
rect 3534 5794 3586 5846
rect 3614 5794 3666 5846
rect 1884 5049 1936 5101
rect 1884 4959 1936 5011
rect 574 4744 626 4796
rect 654 4744 706 4796
rect 944 4744 996 4796
rect 1024 4744 1076 4796
rect 1314 4744 1366 4796
rect 1394 4744 1446 4796
rect 2424 4744 2476 4796
rect 2504 4744 2556 4796
rect 2794 4744 2846 4796
rect 2874 4744 2926 4796
rect 3164 4744 3216 4796
rect 3244 4744 3296 4796
rect 1704 4654 1756 4706
rect 1804 4654 1856 4706
rect 1904 4654 1956 4706
rect 204 4564 256 4616
rect 284 4564 336 4616
rect 574 4564 626 4616
rect 654 4564 706 4616
rect 944 4564 996 4616
rect 1024 4564 1076 4616
rect 1314 4564 1366 4616
rect 1394 4564 1446 4616
rect 1684 4564 1736 4616
rect 1764 4564 1816 4616
rect 574 3514 626 3566
rect 654 3514 706 3566
rect 944 3514 996 3566
rect 1024 3514 1076 3566
rect 1314 3514 1366 3566
rect 1394 3514 1446 3566
rect 2134 4564 2186 4616
rect 2424 4564 2476 4616
rect 2504 4564 2556 4616
rect 2794 4564 2846 4616
rect 2874 4564 2926 4616
rect 3164 4564 3216 4616
rect 3244 4564 3296 4616
rect 3534 4564 3586 4616
rect 3614 4564 3666 4616
rect 2254 3804 2306 3856
rect 2254 3724 2306 3776
rect 2424 3514 2476 3566
rect 2504 3514 2556 3566
rect 2794 3514 2846 3566
rect 2874 3514 2926 3566
rect 3164 3514 3216 3566
rect 3244 3514 3296 3566
rect 204 3394 256 3446
rect 284 3394 336 3446
rect 574 3394 626 3446
rect 654 3394 706 3446
rect 944 3394 996 3446
rect 1024 3394 1076 3446
rect 1314 3394 1366 3446
rect 1394 3394 1446 3446
rect 1684 3394 1736 3446
rect 1764 3394 1816 3446
rect 2054 3394 2106 3446
rect 2134 3394 2186 3446
rect 2424 3394 2476 3446
rect 2504 3394 2556 3446
rect 2794 3394 2846 3446
rect 2874 3394 2926 3446
rect 3164 3394 3216 3446
rect 3244 3394 3296 3446
rect 3534 3394 3586 3446
rect 3614 3394 3666 3446
rect 574 2344 626 2396
rect 654 2344 706 2396
rect 944 2344 996 2396
rect 1024 2344 1076 2396
rect 1314 2344 1366 2396
rect 1394 2344 1446 2396
rect 1684 2344 1736 2396
rect 1764 2344 1816 2396
rect 2054 2344 2106 2396
rect 2134 2344 2186 2396
rect 2424 2344 2476 2396
rect 2504 2344 2556 2396
rect 2794 2344 2846 2396
rect 2874 2344 2926 2396
rect 3164 2344 3216 2396
rect 3244 2344 3296 2396
rect 204 2224 256 2276
rect 284 2224 336 2276
rect 574 2224 626 2276
rect 654 2224 706 2276
rect 944 2224 996 2276
rect 1024 2224 1076 2276
rect 1314 2224 1366 2276
rect 1394 2224 1446 2276
rect 1684 2224 1736 2276
rect 1764 2224 1816 2276
rect 2054 2224 2106 2276
rect 2134 2224 2186 2276
rect 2424 2224 2476 2276
rect 2504 2224 2556 2276
rect 2794 2224 2846 2276
rect 2874 2224 2926 2276
rect 3164 2224 3216 2276
rect 3244 2224 3296 2276
rect 3534 2224 3586 2276
rect 3614 2224 3666 2276
rect 574 1174 626 1226
rect 654 1174 706 1226
rect 944 1174 996 1226
rect 1024 1174 1076 1226
rect 1314 1174 1366 1226
rect 1394 1174 1446 1226
rect 1684 1174 1736 1226
rect 1764 1174 1816 1226
rect 2054 1174 2106 1226
rect 2134 1174 2186 1226
rect 2424 1174 2476 1226
rect 2504 1174 2556 1226
rect 2794 1174 2846 1226
rect 2874 1174 2926 1226
rect 3164 1174 3216 1226
rect 3244 1174 3296 1226
rect 204 1054 256 1106
rect 284 1054 336 1106
rect 574 1054 626 1106
rect 654 1054 706 1106
rect 944 1054 996 1106
rect 1024 1054 1076 1106
rect 1314 1054 1366 1106
rect 1394 1054 1446 1106
rect 1684 1054 1736 1106
rect 1764 1054 1816 1106
rect 2054 1054 2106 1106
rect 2134 1054 2186 1106
rect 2424 1054 2476 1106
rect 2504 1054 2556 1106
rect 2794 1054 2846 1106
rect 2874 1054 2926 1106
rect 3164 1054 3216 1106
rect 3244 1054 3296 1106
rect 3534 1054 3586 1106
rect 3614 1054 3666 1106
rect 574 4 626 56
rect 654 4 706 56
rect 944 4 996 56
rect 1024 4 1076 56
rect 1314 4 1366 56
rect 1394 4 1446 56
rect 1684 4 1736 56
rect 1764 4 1816 56
rect 2054 4 2106 56
rect 2134 4 2186 56
rect 2424 4 2476 56
rect 2504 4 2556 56
rect 2794 4 2846 56
rect 2874 4 2926 56
rect 3164 4 3216 56
rect 3244 4 3296 56
<< metal2 >>
rect 3870 9418 3970 9440
rect 3870 9362 3892 9418
rect 3948 9362 3970 9418
rect 3870 9360 3970 9362
rect 190 9356 3970 9360
rect 190 9304 204 9356
rect 256 9304 284 9356
rect 336 9304 574 9356
rect 626 9304 654 9356
rect 706 9304 944 9356
rect 996 9304 1024 9356
rect 1076 9304 1314 9356
rect 1366 9304 1394 9356
rect 1446 9304 1684 9356
rect 1736 9304 1764 9356
rect 1816 9304 2054 9356
rect 2106 9304 2134 9356
rect 2186 9304 2424 9356
rect 2476 9304 2504 9356
rect 2556 9304 2794 9356
rect 2846 9304 2874 9356
rect 2926 9304 3164 9356
rect 3216 9304 3244 9356
rect 3296 9304 3534 9356
rect 3586 9304 3614 9356
rect 3666 9304 3970 9356
rect 190 9300 3970 9304
rect 3870 9298 3970 9300
rect 3870 9242 3892 9298
rect 3948 9242 3970 9298
rect 3870 9220 3970 9242
rect -60 8368 40 8390
rect -60 8312 -38 8368
rect 18 8312 40 8368
rect -60 8310 40 8312
rect -60 8306 3420 8310
rect -60 8254 574 8306
rect 626 8254 654 8306
rect 706 8254 944 8306
rect 996 8254 1024 8306
rect 1076 8254 1314 8306
rect 1366 8254 1394 8306
rect 1446 8254 1684 8306
rect 1736 8254 1764 8306
rect 1816 8254 2054 8306
rect 2106 8254 2134 8306
rect 2186 8254 2424 8306
rect 2476 8254 2504 8306
rect 2556 8254 2794 8306
rect 2846 8254 2874 8306
rect 2926 8254 3164 8306
rect 3216 8254 3244 8306
rect 3296 8254 3420 8306
rect -60 8250 3420 8254
rect -60 8248 40 8250
rect -60 8192 -38 8248
rect 18 8192 40 8248
rect -60 8170 40 8192
rect 3870 8248 3970 8270
rect 3870 8192 3892 8248
rect 3948 8192 3970 8248
rect 3870 8190 3970 8192
rect 190 8186 3970 8190
rect 190 8134 204 8186
rect 256 8134 284 8186
rect 336 8134 574 8186
rect 626 8134 654 8186
rect 706 8134 944 8186
rect 996 8134 1024 8186
rect 1076 8134 1314 8186
rect 1366 8134 1394 8186
rect 1446 8134 1684 8186
rect 1736 8134 1764 8186
rect 1816 8134 2054 8186
rect 2106 8134 2134 8186
rect 2186 8134 2424 8186
rect 2476 8134 2504 8186
rect 2556 8134 2794 8186
rect 2846 8134 2874 8186
rect 2926 8134 3164 8186
rect 3216 8134 3244 8186
rect 3296 8134 3534 8186
rect 3586 8134 3614 8186
rect 3666 8134 3970 8186
rect 190 8130 3970 8134
rect 3870 8128 3970 8130
rect 3870 8072 3892 8128
rect 3948 8072 3970 8128
rect 3870 8050 3970 8072
rect -60 7198 40 7220
rect -60 7142 -38 7198
rect 18 7142 40 7198
rect -60 7140 40 7142
rect -60 7136 3420 7140
rect -60 7084 574 7136
rect 626 7084 654 7136
rect 706 7084 944 7136
rect 996 7084 1024 7136
rect 1076 7084 1314 7136
rect 1366 7084 1394 7136
rect 1446 7084 1684 7136
rect 1736 7084 1764 7136
rect 1816 7084 2054 7136
rect 2106 7084 2134 7136
rect 2186 7084 2424 7136
rect 2476 7084 2504 7136
rect 2556 7084 2794 7136
rect 2846 7084 2874 7136
rect 2926 7084 3164 7136
rect 3216 7084 3244 7136
rect 3296 7084 3420 7136
rect -60 7080 3420 7084
rect -60 7078 40 7080
rect -60 7022 -38 7078
rect 18 7022 40 7078
rect -60 7000 40 7022
rect 3870 7078 3970 7100
rect 3870 7022 3892 7078
rect 3948 7022 3970 7078
rect 3870 7020 3970 7022
rect 190 7016 3970 7020
rect 190 6964 204 7016
rect 256 6964 284 7016
rect 336 6964 574 7016
rect 626 6964 654 7016
rect 706 6964 944 7016
rect 996 6964 1024 7016
rect 1076 6964 1314 7016
rect 1366 6964 1394 7016
rect 1446 6964 1684 7016
rect 1736 6964 1764 7016
rect 1816 6964 2054 7016
rect 2106 6964 2134 7016
rect 2186 6964 2424 7016
rect 2476 6964 2504 7016
rect 2556 6964 2794 7016
rect 2846 6964 2874 7016
rect 2926 6964 3164 7016
rect 3216 6964 3244 7016
rect 3296 6964 3534 7016
rect 3586 6964 3614 7016
rect 3666 6964 3970 7016
rect 190 6960 3970 6964
rect 3870 6958 3970 6960
rect 3870 6902 3892 6958
rect 3948 6902 3970 6958
rect 3870 6880 3970 6902
rect -60 6028 40 6050
rect -60 5972 -38 6028
rect 18 5972 40 6028
rect -60 5970 40 5972
rect 3870 5988 3970 6010
rect -60 5966 3420 5970
rect -60 5914 574 5966
rect 626 5914 654 5966
rect 706 5914 944 5966
rect 996 5914 1024 5966
rect 1076 5914 1314 5966
rect 1366 5914 1394 5966
rect 1446 5914 1684 5966
rect 1736 5914 1764 5966
rect 1816 5914 2054 5966
rect 2106 5914 2134 5966
rect 2186 5914 2424 5966
rect 2476 5914 2504 5966
rect 2556 5914 2794 5966
rect 2846 5914 2874 5966
rect 2926 5914 3164 5966
rect 3216 5914 3244 5966
rect 3296 5914 3420 5966
rect -60 5910 3420 5914
rect 3870 5932 3892 5988
rect 3948 5932 3970 5988
rect -60 5908 40 5910
rect -60 5852 -38 5908
rect 18 5852 40 5908
rect -60 5830 40 5852
rect 3870 5868 3970 5932
rect 3870 5850 3892 5868
rect 190 5846 3892 5850
rect 190 5794 204 5846
rect 256 5794 284 5846
rect 336 5794 574 5846
rect 626 5794 654 5846
rect 706 5794 944 5846
rect 996 5794 1024 5846
rect 1076 5794 1314 5846
rect 1366 5794 1394 5846
rect 1446 5794 1684 5846
rect 1736 5794 1764 5846
rect 1816 5794 2054 5846
rect 2106 5794 2134 5846
rect 2186 5794 2424 5846
rect 2476 5794 2504 5846
rect 2556 5794 2794 5846
rect 2846 5794 2874 5846
rect 2926 5794 3164 5846
rect 3216 5794 3244 5846
rect 3296 5794 3534 5846
rect 3586 5794 3614 5846
rect 3666 5812 3892 5846
rect 3948 5812 3970 5868
rect 3666 5794 3970 5812
rect 190 5790 3970 5794
rect 1880 5101 1940 5120
rect 1880 5049 1884 5101
rect 1936 5049 1940 5101
rect 1880 5011 1940 5049
rect -60 4938 40 4960
rect -60 4882 -38 4938
rect 18 4882 40 4938
rect -60 4818 40 4882
rect -60 4762 -38 4818
rect 18 4800 40 4818
rect 1880 4959 1884 5011
rect 1936 4959 1940 5011
rect 1880 4800 1940 4959
rect 18 4796 3420 4800
rect 18 4762 574 4796
rect -60 4744 574 4762
rect 626 4744 654 4796
rect 706 4744 944 4796
rect 996 4744 1024 4796
rect 1076 4744 1314 4796
rect 1366 4744 1394 4796
rect 1446 4744 2424 4796
rect 2476 4744 2504 4796
rect 2556 4744 2794 4796
rect 2846 4744 2874 4796
rect 2926 4744 3164 4796
rect 3216 4744 3244 4796
rect 3296 4744 3420 4796
rect -60 4740 3420 4744
rect -240 4710 -140 4730
rect -240 4708 2020 4710
rect -240 4652 -218 4708
rect -162 4706 2020 4708
rect -162 4654 1704 4706
rect 1756 4654 1804 4706
rect 1856 4654 1904 4706
rect 1956 4654 2020 4706
rect -162 4652 2020 4654
rect -240 4650 2020 4652
rect 3870 4678 3970 4700
rect -240 4630 -140 4650
rect 3870 4622 3892 4678
rect 3948 4622 3970 4678
rect 3870 4620 3970 4622
rect 190 4616 3970 4620
rect 190 4564 204 4616
rect 256 4564 284 4616
rect 336 4564 574 4616
rect 626 4564 654 4616
rect 706 4564 944 4616
rect 996 4564 1024 4616
rect 1076 4564 1314 4616
rect 1366 4564 1394 4616
rect 1446 4564 1684 4616
rect 1736 4564 1764 4616
rect 1816 4564 2134 4616
rect 2186 4564 2424 4616
rect 2476 4564 2504 4616
rect 2556 4564 2794 4616
rect 2846 4564 2874 4616
rect 2926 4564 3164 4616
rect 3216 4564 3244 4616
rect 3296 4564 3534 4616
rect 3586 4564 3614 4616
rect 3666 4564 3970 4616
rect 190 4560 3970 4564
rect 3870 4558 3970 4560
rect 3870 4502 3892 4558
rect 3948 4502 3970 4558
rect 3870 4480 3970 4502
rect 2250 3856 2310 3880
rect 2250 3804 2254 3856
rect 2306 3804 2310 3856
rect 2250 3776 2310 3804
rect 2250 3724 2254 3776
rect 2306 3724 2310 3776
rect -60 3628 40 3650
rect -60 3572 -38 3628
rect 18 3572 40 3628
rect -60 3570 40 3572
rect 2250 3570 2310 3724
rect -60 3566 3420 3570
rect -60 3514 574 3566
rect 626 3514 654 3566
rect 706 3514 944 3566
rect 996 3514 1024 3566
rect 1076 3514 1314 3566
rect 1366 3514 1394 3566
rect 1446 3514 2424 3566
rect 2476 3514 2504 3566
rect 2556 3514 2794 3566
rect 2846 3514 2874 3566
rect 2926 3514 3164 3566
rect 3216 3514 3244 3566
rect 3296 3514 3420 3566
rect -60 3510 3420 3514
rect -60 3508 40 3510
rect -60 3452 -38 3508
rect 18 3452 40 3508
rect -60 3430 40 3452
rect 3870 3508 3970 3530
rect 3870 3452 3892 3508
rect 3948 3452 3970 3508
rect 3870 3450 3970 3452
rect 190 3446 3970 3450
rect 190 3394 204 3446
rect 256 3394 284 3446
rect 336 3394 574 3446
rect 626 3394 654 3446
rect 706 3394 944 3446
rect 996 3394 1024 3446
rect 1076 3394 1314 3446
rect 1366 3394 1394 3446
rect 1446 3394 1684 3446
rect 1736 3394 1764 3446
rect 1816 3394 2054 3446
rect 2106 3394 2134 3446
rect 2186 3394 2424 3446
rect 2476 3394 2504 3446
rect 2556 3394 2794 3446
rect 2846 3394 2874 3446
rect 2926 3394 3164 3446
rect 3216 3394 3244 3446
rect 3296 3394 3534 3446
rect 3586 3394 3614 3446
rect 3666 3394 3970 3446
rect 190 3390 3970 3394
rect 3870 3388 3970 3390
rect 3870 3332 3892 3388
rect 3948 3332 3970 3388
rect 3870 3310 3970 3332
rect -60 2458 40 2480
rect -60 2402 -38 2458
rect 18 2402 40 2458
rect -60 2400 40 2402
rect -60 2396 3420 2400
rect -60 2344 574 2396
rect 626 2344 654 2396
rect 706 2344 944 2396
rect 996 2344 1024 2396
rect 1076 2344 1314 2396
rect 1366 2344 1394 2396
rect 1446 2344 1684 2396
rect 1736 2344 1764 2396
rect 1816 2344 2054 2396
rect 2106 2344 2134 2396
rect 2186 2344 2424 2396
rect 2476 2344 2504 2396
rect 2556 2344 2794 2396
rect 2846 2344 2874 2396
rect 2926 2344 3164 2396
rect 3216 2344 3244 2396
rect 3296 2344 3420 2396
rect -60 2340 3420 2344
rect -60 2338 40 2340
rect -60 2282 -38 2338
rect 18 2282 40 2338
rect -60 2260 40 2282
rect 3870 2338 3970 2360
rect 3870 2282 3892 2338
rect 3948 2282 3970 2338
rect 3870 2280 3970 2282
rect 190 2276 3970 2280
rect 190 2224 204 2276
rect 256 2224 284 2276
rect 336 2224 574 2276
rect 626 2224 654 2276
rect 706 2224 944 2276
rect 996 2224 1024 2276
rect 1076 2224 1314 2276
rect 1366 2224 1394 2276
rect 1446 2224 1684 2276
rect 1736 2224 1764 2276
rect 1816 2224 2054 2276
rect 2106 2224 2134 2276
rect 2186 2224 2424 2276
rect 2476 2224 2504 2276
rect 2556 2224 2794 2276
rect 2846 2224 2874 2276
rect 2926 2224 3164 2276
rect 3216 2224 3244 2276
rect 3296 2224 3534 2276
rect 3586 2224 3614 2276
rect 3666 2224 3970 2276
rect 190 2220 3970 2224
rect 3870 2218 3970 2220
rect 3870 2162 3892 2218
rect 3948 2162 3970 2218
rect 3870 2140 3970 2162
rect -60 1288 40 1310
rect -60 1232 -38 1288
rect 18 1232 40 1288
rect -60 1230 40 1232
rect -60 1226 3420 1230
rect -60 1174 574 1226
rect 626 1174 654 1226
rect 706 1174 944 1226
rect 996 1174 1024 1226
rect 1076 1174 1314 1226
rect 1366 1174 1394 1226
rect 1446 1174 1684 1226
rect 1736 1174 1764 1226
rect 1816 1174 2054 1226
rect 2106 1174 2134 1226
rect 2186 1174 2424 1226
rect 2476 1174 2504 1226
rect 2556 1174 2794 1226
rect 2846 1174 2874 1226
rect 2926 1174 3164 1226
rect 3216 1174 3244 1226
rect 3296 1174 3420 1226
rect -60 1170 3420 1174
rect -60 1168 40 1170
rect -60 1112 -38 1168
rect 18 1112 40 1168
rect -60 1090 40 1112
rect 3870 1168 3970 1190
rect 3870 1112 3892 1168
rect 3948 1112 3970 1168
rect 3870 1110 3970 1112
rect 190 1106 3970 1110
rect 190 1054 204 1106
rect 256 1054 284 1106
rect 336 1054 574 1106
rect 626 1054 654 1106
rect 706 1054 944 1106
rect 996 1054 1024 1106
rect 1076 1054 1314 1106
rect 1366 1054 1394 1106
rect 1446 1054 1684 1106
rect 1736 1054 1764 1106
rect 1816 1054 2054 1106
rect 2106 1054 2134 1106
rect 2186 1054 2424 1106
rect 2476 1054 2504 1106
rect 2556 1054 2794 1106
rect 2846 1054 2874 1106
rect 2926 1054 3164 1106
rect 3216 1054 3244 1106
rect 3296 1054 3534 1106
rect 3586 1054 3614 1106
rect 3666 1054 3970 1106
rect 190 1050 3970 1054
rect 3870 1048 3970 1050
rect 3870 992 3892 1048
rect 3948 992 3970 1048
rect 3870 970 3970 992
rect -60 118 40 140
rect -60 62 -38 118
rect 18 62 40 118
rect -60 60 40 62
rect -60 56 3420 60
rect -60 4 574 56
rect 626 4 654 56
rect 706 4 944 56
rect 996 4 1024 56
rect 1076 4 1314 56
rect 1366 4 1394 56
rect 1446 4 1684 56
rect 1736 4 1764 56
rect 1816 4 2054 56
rect 2106 4 2134 56
rect 2186 4 2424 56
rect 2476 4 2504 56
rect 2556 4 2794 56
rect 2846 4 2874 56
rect 2926 4 3164 56
rect 3216 4 3244 56
rect 3296 4 3420 56
rect -60 0 3420 4
rect -60 -2 40 0
rect -60 -58 -38 -2
rect 18 -58 40 -2
rect -60 -80 40 -58
<< via2 >>
rect 3892 9362 3948 9418
rect 3892 9242 3948 9298
rect -38 8312 18 8368
rect -38 8192 18 8248
rect 3892 8192 3948 8248
rect 3892 8072 3948 8128
rect -38 7142 18 7198
rect -38 7022 18 7078
rect 3892 7022 3948 7078
rect 3892 6902 3948 6958
rect -38 5972 18 6028
rect 3892 5932 3948 5988
rect -38 5852 18 5908
rect 3892 5812 3948 5868
rect -38 4882 18 4938
rect -38 4762 18 4818
rect -218 4652 -162 4708
rect 3892 4622 3948 4678
rect 3892 4502 3948 4558
rect -38 3572 18 3628
rect -38 3452 18 3508
rect 3892 3452 3948 3508
rect 3892 3332 3948 3388
rect -38 2402 18 2458
rect -38 2282 18 2338
rect 3892 2282 3948 2338
rect 3892 2162 3948 2218
rect -38 1232 18 1288
rect -38 1112 18 1168
rect 3892 1112 3948 1168
rect 3892 992 3948 1048
rect -38 62 18 118
rect -38 -58 18 -2
<< metal3 >>
rect -60 8368 40 9820
rect -60 8312 -38 8368
rect 18 8312 40 8368
rect -60 8248 40 8312
rect -60 8192 -38 8248
rect 18 8192 40 8248
rect -60 7198 40 8192
rect -60 7142 -38 7198
rect 18 7142 40 7198
rect -60 7078 40 7142
rect -60 7022 -38 7078
rect 18 7022 40 7078
rect -60 6028 40 7022
rect -60 5972 -38 6028
rect 18 5972 40 6028
rect -60 5908 40 5972
rect -60 5852 -38 5908
rect 18 5852 40 5908
rect -60 4938 40 5852
rect -60 4882 -38 4938
rect 18 4882 40 4938
rect -60 4818 40 4882
rect -60 4762 -38 4818
rect 18 4762 40 4818
rect -240 4708 -140 4730
rect -240 4652 -218 4708
rect -162 4652 -140 4708
rect -240 4630 -140 4652
rect -60 3628 40 4762
rect -60 3572 -38 3628
rect 18 3572 40 3628
rect -60 3508 40 3572
rect -60 3452 -38 3508
rect 18 3452 40 3508
rect -60 2458 40 3452
rect -60 2402 -38 2458
rect 18 2402 40 2458
rect -60 2338 40 2402
rect -60 2282 -38 2338
rect 18 2282 40 2338
rect -60 1288 40 2282
rect -60 1232 -38 1288
rect 18 1232 40 1288
rect -60 1168 40 1232
rect -60 1112 -38 1168
rect 18 1112 40 1168
rect -60 118 40 1112
rect 3870 9418 3970 9697
rect 3870 9362 3892 9418
rect 3948 9362 3970 9418
rect 3870 9298 3970 9362
rect 3870 9242 3892 9298
rect 3948 9242 3970 9298
rect 3870 8248 3970 9242
rect 3870 8192 3892 8248
rect 3948 8192 3970 8248
rect 3870 8128 3970 8192
rect 3870 8072 3892 8128
rect 3948 8072 3970 8128
rect 3870 7078 3970 8072
rect 3870 7022 3892 7078
rect 3948 7022 3970 7078
rect 3870 6958 3970 7022
rect 3870 6902 3892 6958
rect 3948 6902 3970 6958
rect 3870 5988 3970 6902
rect 3870 5932 3892 5988
rect 3948 5932 3970 5988
rect 3870 5868 3970 5932
rect 3870 5812 3892 5868
rect 3948 5812 3970 5868
rect 3870 4678 3970 5812
rect 3870 4622 3892 4678
rect 3948 4622 3970 4678
rect 3870 4558 3970 4622
rect 3870 4502 3892 4558
rect 3948 4502 3970 4558
rect 3870 3508 3970 4502
rect 3870 3452 3892 3508
rect 3948 3452 3970 3508
rect 3870 3388 3970 3452
rect 3870 3332 3892 3388
rect 3948 3332 3970 3388
rect 3870 2338 3970 3332
rect 3870 2282 3892 2338
rect 3948 2282 3970 2338
rect 3870 2218 3970 2282
rect 3870 2162 3892 2218
rect 3948 2162 3970 2218
rect 3870 1168 3970 2162
rect 3870 1112 3892 1168
rect 3948 1112 3970 1168
rect 3870 1048 3970 1112
rect 3870 992 3892 1048
rect 3948 992 3970 1048
rect 3870 970 3970 992
rect -60 62 -38 118
rect 18 62 40 118
rect -60 -2 40 62
rect -60 -58 -38 -2
rect 18 -58 40 -2
rect -60 -80 40 -58
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_0
timestamp 1757161594
transform 0 1 3638 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_1
timestamp 1757161594
transform 0 1 2528 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_2
timestamp 1757161594
transform 0 1 2898 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_3
timestamp 1757161594
transform 0 1 1048 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_4
timestamp 1757161594
transform 0 1 678 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_5
timestamp 1757161594
transform 0 1 308 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_6
timestamp 1757161594
transform 0 1 1418 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_7
timestamp 1757161594
transform 0 1 1788 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_8
timestamp 1757161594
transform 0 1 2158 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_9
timestamp 1757161594
transform 0 1 3268 1 0 554
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_10
timestamp 1757161594
transform 0 1 3638 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_11
timestamp 1757161594
transform 0 1 3268 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_12
timestamp 1757161594
transform 0 1 2898 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_13
timestamp 1757161594
transform 0 1 2528 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_14
timestamp 1757161594
transform 0 1 2158 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_15
timestamp 1757161594
transform 0 1 1788 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_16
timestamp 1757161594
transform 0 1 1418 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_17
timestamp 1757161594
transform 0 1 1048 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_18
timestamp 1757161594
transform 0 1 678 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_19
timestamp 1757161594
transform 0 1 308 1 0 1724
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_20
timestamp 1757161594
transform 0 1 1048 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_21
timestamp 1757161594
transform 0 1 678 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_22
timestamp 1757161594
transform 0 1 308 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_23
timestamp 1757161594
transform 0 1 2158 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_24
timestamp 1757161594
transform 0 1 1788 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_25
timestamp 1757161594
transform 0 1 1418 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_26
timestamp 1757161594
transform 0 1 3638 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_27
timestamp 1757161594
transform 0 1 3268 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_28
timestamp 1757161594
transform 0 1 2898 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_29
timestamp 1757161594
transform 0 1 2528 1 0 2894
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_30
timestamp 1757161594
transform 0 1 3638 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_31
timestamp 1757161594
transform 0 1 3268 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_32
timestamp 1757161594
transform 0 1 2898 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_33
timestamp 1757161594
transform 0 1 2528 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_34
timestamp 1757161594
transform 0 1 2158 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_35
timestamp 1757161594
transform 0 1 1788 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_36
timestamp 1757161594
transform 0 1 1418 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_37
timestamp 1757161594
transform 0 1 1048 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_38
timestamp 1757161594
transform 0 1 678 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_39
timestamp 1757161594
transform 0 1 308 1 0 4064
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_40
timestamp 1757161594
transform 0 1 1048 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_41
timestamp 1757161594
transform 0 1 678 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_42
timestamp 1757161594
transform 0 1 308 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_43
timestamp 1757161594
transform 0 1 2158 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_44
timestamp 1757161594
transform 0 1 1788 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_45
timestamp 1757161594
transform 0 1 1418 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_46
timestamp 1757161594
transform 0 1 3638 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_47
timestamp 1757161594
transform 0 1 3268 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_48
timestamp 1757161594
transform 0 1 2898 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_49
timestamp 1757161594
transform 0 1 2528 1 0 5294
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_50
timestamp 1757161594
transform 0 1 3638 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_51
timestamp 1757161594
transform 0 1 3268 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_52
timestamp 1757161594
transform 0 1 2898 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_53
timestamp 1757161594
transform 0 1 2528 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_54
timestamp 1757161594
transform 0 1 2158 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_55
timestamp 1757161594
transform 0 1 1788 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_56
timestamp 1757161594
transform 0 1 1418 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_57
timestamp 1757161594
transform 0 1 1048 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_58
timestamp 1757161594
transform 0 1 678 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_59
timestamp 1757161594
transform 0 1 308 1 0 6464
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_60
timestamp 1757161594
transform 0 1 1048 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_61
timestamp 1757161594
transform 0 1 678 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_62
timestamp 1757161594
transform 0 1 308 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_63
timestamp 1757161594
transform 0 1 2158 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_64
timestamp 1757161594
transform 0 1 1788 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_65
timestamp 1757161594
transform 0 1 1418 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_66
timestamp 1757161594
transform 0 1 3638 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_67
timestamp 1757161594
transform 0 1 3268 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_68
timestamp 1757161594
transform 0 1 2898 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_69
timestamp 1757161594
transform 0 1 2528 1 0 8804
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_70
timestamp 1757161594
transform 0 1 1048 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_71
timestamp 1757161594
transform 0 1 678 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_72
timestamp 1757161594
transform 0 1 308 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_73
timestamp 1757161594
transform 0 1 2158 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_74
timestamp 1757161594
transform 0 1 1788 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_75
timestamp 1757161594
transform 0 1 1418 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_76
timestamp 1757161594
transform 0 1 3638 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_77
timestamp 1757161594
transform 0 1 3268 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_78
timestamp 1757161594
transform 0 1 2898 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_KVZN99  sky130_fd_pr__pfet_01v8_lvt_KVZN99_79
timestamp 1757161594
transform 0 1 2528 1 0 7634
box -594 -198 594 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_0
timestamp 1757161594
transform 0 1 1048 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_1
timestamp 1757161594
transform 0 1 308 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_2
timestamp 1757161594
transform 0 1 678 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_3
timestamp 1757161594
transform 0 1 2158 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_4
timestamp 1757161594
transform 0 1 1418 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_5
timestamp 1757161594
transform 0 1 1788 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_6
timestamp 1757161594
transform 0 1 2898 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_7
timestamp 1757161594
transform 0 1 3638 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_8
timestamp 1757161594
transform 0 1 2528 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_9
timestamp 1757161594
transform 0 1 3268 1 0 -166
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_10
timestamp 1757161594
transform 0 1 1048 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_11
timestamp 1757161594
transform 0 1 678 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_12
timestamp 1757161594
transform 0 1 308 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_13
timestamp 1757161594
transform 0 1 2158 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_14
timestamp 1757161594
transform 0 1 1418 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_15
timestamp 1757161594
transform 0 1 1788 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_16
timestamp 1757161594
transform 0 1 3638 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_17
timestamp 1757161594
transform 0 1 2898 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_18
timestamp 1757161594
transform 0 1 3268 1 0 9524
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_lvt_MTZNSY  sky130_fd_pr__pfet_01v8_lvt_MTZNSY_19
timestamp 1757161594
transform 0 1 2528 1 0 9524
box -144 -198 144 164
<< labels >>
flabel metal3 s -60 9720 40 9820 0 FreeSans 1172 0 0 0 Vb
port 0 nsew
<< end >>
