magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -386 -369 386 369
<< nmoslvt >>
rect -200 -231 200 169
<< ndiff >>
rect -258 156 -200 169
rect -258 122 -246 156
rect -212 122 -200 156
rect -258 88 -200 122
rect -258 54 -246 88
rect -212 54 -200 88
rect -258 20 -200 54
rect -258 -14 -246 20
rect -212 -14 -200 20
rect -258 -48 -200 -14
rect -258 -82 -246 -48
rect -212 -82 -200 -48
rect -258 -116 -200 -82
rect -258 -150 -246 -116
rect -212 -150 -200 -116
rect -258 -184 -200 -150
rect -258 -218 -246 -184
rect -212 -218 -200 -184
rect -258 -231 -200 -218
rect 200 156 258 169
rect 200 122 212 156
rect 246 122 258 156
rect 200 88 258 122
rect 200 54 212 88
rect 246 54 258 88
rect 200 20 258 54
rect 200 -14 212 20
rect 246 -14 258 20
rect 200 -48 258 -14
rect 200 -82 212 -48
rect 246 -82 258 -48
rect 200 -116 258 -82
rect 200 -150 212 -116
rect 246 -150 258 -116
rect 200 -184 258 -150
rect 200 -218 212 -184
rect 246 -218 258 -184
rect 200 -231 258 -218
<< ndiffc >>
rect -246 122 -212 156
rect -246 54 -212 88
rect -246 -14 -212 20
rect -246 -82 -212 -48
rect -246 -150 -212 -116
rect -246 -218 -212 -184
rect 212 122 246 156
rect 212 54 246 88
rect 212 -14 246 20
rect 212 -82 246 -48
rect 212 -150 246 -116
rect 212 -218 246 -184
<< psubdiff >>
rect -360 309 360 343
rect -360 -309 -326 309
rect 326 -309 360 309
rect -360 -343 -255 -309
rect -221 -343 -187 -309
rect -153 -343 -119 -309
rect -85 -343 -51 -309
rect -17 -343 17 -309
rect 51 -343 85 -309
rect 119 -343 153 -309
rect 187 -343 221 -309
rect 255 -343 360 -309
<< psubdiffcont >>
rect -255 -343 -221 -309
rect -187 -343 -153 -309
rect -119 -343 -85 -309
rect -51 -343 -17 -309
rect 17 -343 51 -309
rect 85 -343 119 -309
rect 153 -343 187 -309
rect 221 -343 255 -309
<< poly >>
rect -200 241 200 257
rect -200 207 -153 241
rect -119 207 -85 241
rect -51 207 -17 241
rect 17 207 51 241
rect 85 207 119 241
rect 153 207 200 241
rect -200 169 200 207
rect -200 -257 200 -231
<< polycont >>
rect -153 207 -119 241
rect -85 207 -51 241
rect -17 207 17 241
rect 51 207 85 241
rect 119 207 153 241
<< locali >>
rect -360 309 360 343
rect -360 -309 -326 309
rect -200 207 -161 241
rect -119 207 -89 241
rect -51 207 -17 241
rect 17 207 51 241
rect 89 207 119 241
rect 161 207 200 241
rect -246 156 -212 173
rect -246 88 -212 96
rect -246 20 -212 24
rect -246 -86 -212 -82
rect -246 -158 -212 -150
rect -246 -235 -212 -218
rect 212 156 246 173
rect 212 88 246 96
rect 212 20 246 24
rect 212 -86 246 -82
rect 212 -158 246 -150
rect 212 -235 246 -218
rect 326 -309 360 309
rect -360 -343 -255 -309
rect -221 -343 -187 -309
rect -153 -343 -119 -309
rect -85 -343 -51 -309
rect -17 -343 17 -309
rect 51 -343 85 -309
rect 119 -343 153 -309
rect 187 -343 221 -309
rect 255 -343 360 -309
<< viali >>
rect -161 207 -153 241
rect -153 207 -127 241
rect -89 207 -85 241
rect -85 207 -55 241
rect -17 207 17 241
rect 55 207 85 241
rect 85 207 89 241
rect 127 207 153 241
rect 153 207 161 241
rect -246 122 -212 130
rect -246 96 -212 122
rect -246 54 -212 58
rect -246 24 -212 54
rect -246 -48 -212 -14
rect -246 -116 -212 -86
rect -246 -120 -212 -116
rect -246 -184 -212 -158
rect -246 -192 -212 -184
rect 212 122 246 130
rect 212 96 246 122
rect 212 54 246 58
rect 212 24 246 54
rect 212 -48 246 -14
rect 212 -116 246 -86
rect 212 -120 246 -116
rect 212 -184 246 -158
rect 212 -192 246 -184
<< metal1 >>
rect -196 241 196 247
rect -196 207 -161 241
rect -127 207 -89 241
rect -55 207 -17 241
rect 17 207 55 241
rect 89 207 127 241
rect 161 207 196 241
rect -196 201 196 207
rect -252 130 -206 169
rect -252 96 -246 130
rect -212 96 -206 130
rect -252 58 -206 96
rect -252 24 -246 58
rect -212 24 -206 58
rect -252 -14 -206 24
rect -252 -48 -246 -14
rect -212 -48 -206 -14
rect -252 -86 -206 -48
rect -252 -120 -246 -86
rect -212 -120 -206 -86
rect -252 -158 -206 -120
rect -252 -192 -246 -158
rect -212 -192 -206 -158
rect -252 -231 -206 -192
rect 206 130 252 169
rect 206 96 212 130
rect 246 96 252 130
rect 206 58 252 96
rect 206 24 212 58
rect 246 24 252 58
rect 206 -14 252 24
rect 206 -48 212 -14
rect 246 -48 252 -14
rect 206 -86 252 -48
rect 206 -120 212 -86
rect 246 -120 252 -86
rect 206 -158 252 -120
rect 206 -192 212 -158
rect 246 -192 252 -158
rect 206 -231 252 -192
<< properties >>
string FIXED_BBOX -343 -326 343 326
<< end >>
