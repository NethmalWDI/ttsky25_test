magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -194 -598 194 564
<< pmoslvt >>
rect -100 -536 100 464
<< pdiff >>
rect -158 423 -100 464
rect -158 389 -146 423
rect -112 389 -100 423
rect -158 355 -100 389
rect -158 321 -146 355
rect -112 321 -100 355
rect -158 287 -100 321
rect -158 253 -146 287
rect -112 253 -100 287
rect -158 219 -100 253
rect -158 185 -146 219
rect -112 185 -100 219
rect -158 151 -100 185
rect -158 117 -146 151
rect -112 117 -100 151
rect -158 83 -100 117
rect -158 49 -146 83
rect -112 49 -100 83
rect -158 15 -100 49
rect -158 -19 -146 15
rect -112 -19 -100 15
rect -158 -53 -100 -19
rect -158 -87 -146 -53
rect -112 -87 -100 -53
rect -158 -121 -100 -87
rect -158 -155 -146 -121
rect -112 -155 -100 -121
rect -158 -189 -100 -155
rect -158 -223 -146 -189
rect -112 -223 -100 -189
rect -158 -257 -100 -223
rect -158 -291 -146 -257
rect -112 -291 -100 -257
rect -158 -325 -100 -291
rect -158 -359 -146 -325
rect -112 -359 -100 -325
rect -158 -393 -100 -359
rect -158 -427 -146 -393
rect -112 -427 -100 -393
rect -158 -461 -100 -427
rect -158 -495 -146 -461
rect -112 -495 -100 -461
rect -158 -536 -100 -495
rect 100 423 158 464
rect 100 389 112 423
rect 146 389 158 423
rect 100 355 158 389
rect 100 321 112 355
rect 146 321 158 355
rect 100 287 158 321
rect 100 253 112 287
rect 146 253 158 287
rect 100 219 158 253
rect 100 185 112 219
rect 146 185 158 219
rect 100 151 158 185
rect 100 117 112 151
rect 146 117 158 151
rect 100 83 158 117
rect 100 49 112 83
rect 146 49 158 83
rect 100 15 158 49
rect 100 -19 112 15
rect 146 -19 158 15
rect 100 -53 158 -19
rect 100 -87 112 -53
rect 146 -87 158 -53
rect 100 -121 158 -87
rect 100 -155 112 -121
rect 146 -155 158 -121
rect 100 -189 158 -155
rect 100 -223 112 -189
rect 146 -223 158 -189
rect 100 -257 158 -223
rect 100 -291 112 -257
rect 146 -291 158 -257
rect 100 -325 158 -291
rect 100 -359 112 -325
rect 146 -359 158 -325
rect 100 -393 158 -359
rect 100 -427 112 -393
rect 146 -427 158 -393
rect 100 -461 158 -427
rect 100 -495 112 -461
rect 146 -495 158 -461
rect 100 -536 158 -495
<< pdiffc >>
rect -146 389 -112 423
rect -146 321 -112 355
rect -146 253 -112 287
rect -146 185 -112 219
rect -146 117 -112 151
rect -146 49 -112 83
rect -146 -19 -112 15
rect -146 -87 -112 -53
rect -146 -155 -112 -121
rect -146 -223 -112 -189
rect -146 -291 -112 -257
rect -146 -359 -112 -325
rect -146 -427 -112 -393
rect -146 -495 -112 -461
rect 112 389 146 423
rect 112 321 146 355
rect 112 253 146 287
rect 112 185 146 219
rect 112 117 146 151
rect 112 49 146 83
rect 112 -19 146 15
rect 112 -87 146 -53
rect 112 -155 146 -121
rect 112 -223 146 -189
rect 112 -291 146 -257
rect 112 -359 146 -325
rect 112 -427 146 -393
rect 112 -495 146 -461
<< poly >>
rect -100 545 100 561
rect -100 511 -51 545
rect -17 511 17 545
rect 51 511 100 545
rect -100 464 100 511
rect -100 -562 100 -536
<< polycont >>
rect -51 511 -17 545
rect 17 511 51 545
<< locali >>
rect -100 511 -53 545
rect -17 511 17 545
rect 53 511 100 545
rect -146 449 -112 468
rect -146 377 -112 389
rect -146 305 -112 321
rect -146 233 -112 253
rect -146 161 -112 185
rect -146 89 -112 117
rect -146 17 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -89
rect -146 -189 -112 -161
rect -146 -257 -112 -233
rect -146 -325 -112 -305
rect -146 -393 -112 -377
rect -146 -461 -112 -449
rect -146 -540 -112 -521
rect 112 449 146 468
rect 112 377 146 389
rect 112 305 146 321
rect 112 233 146 253
rect 112 161 146 185
rect 112 89 146 117
rect 112 17 146 49
rect 112 -53 146 -19
rect 112 -121 146 -89
rect 112 -189 146 -161
rect 112 -257 146 -233
rect 112 -325 146 -305
rect 112 -393 146 -377
rect 112 -461 146 -449
rect 112 -540 146 -521
<< viali >>
rect -53 511 -51 545
rect -51 511 -19 545
rect 19 511 51 545
rect 51 511 53 545
rect -146 423 -112 449
rect -146 415 -112 423
rect -146 355 -112 377
rect -146 343 -112 355
rect -146 287 -112 305
rect -146 271 -112 287
rect -146 219 -112 233
rect -146 199 -112 219
rect -146 151 -112 161
rect -146 127 -112 151
rect -146 83 -112 89
rect -146 55 -112 83
rect -146 15 -112 17
rect -146 -17 -112 15
rect -146 -87 -112 -55
rect -146 -89 -112 -87
rect -146 -155 -112 -127
rect -146 -161 -112 -155
rect -146 -223 -112 -199
rect -146 -233 -112 -223
rect -146 -291 -112 -271
rect -146 -305 -112 -291
rect -146 -359 -112 -343
rect -146 -377 -112 -359
rect -146 -427 -112 -415
rect -146 -449 -112 -427
rect -146 -495 -112 -487
rect -146 -521 -112 -495
rect 112 423 146 449
rect 112 415 146 423
rect 112 355 146 377
rect 112 343 146 355
rect 112 287 146 305
rect 112 271 146 287
rect 112 219 146 233
rect 112 199 146 219
rect 112 151 146 161
rect 112 127 146 151
rect 112 83 146 89
rect 112 55 146 83
rect 112 15 146 17
rect 112 -17 146 15
rect 112 -87 146 -55
rect 112 -89 146 -87
rect 112 -155 146 -127
rect 112 -161 146 -155
rect 112 -223 146 -199
rect 112 -233 146 -223
rect 112 -291 146 -271
rect 112 -305 146 -291
rect 112 -359 146 -343
rect 112 -377 146 -359
rect 112 -427 146 -415
rect 112 -449 146 -427
rect 112 -495 146 -487
rect 112 -521 146 -495
<< metal1 >>
rect -96 545 96 551
rect -96 511 -53 545
rect -19 511 19 545
rect 53 511 96 545
rect -96 505 96 511
rect -152 449 -106 464
rect -152 415 -146 449
rect -112 415 -106 449
rect -152 377 -106 415
rect -152 343 -146 377
rect -112 343 -106 377
rect -152 305 -106 343
rect -152 271 -146 305
rect -112 271 -106 305
rect -152 233 -106 271
rect -152 199 -146 233
rect -112 199 -106 233
rect -152 161 -106 199
rect -152 127 -146 161
rect -112 127 -106 161
rect -152 89 -106 127
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -127 -106 -89
rect -152 -161 -146 -127
rect -112 -161 -106 -127
rect -152 -199 -106 -161
rect -152 -233 -146 -199
rect -112 -233 -106 -199
rect -152 -271 -106 -233
rect -152 -305 -146 -271
rect -112 -305 -106 -271
rect -152 -343 -106 -305
rect -152 -377 -146 -343
rect -112 -377 -106 -343
rect -152 -415 -106 -377
rect -152 -449 -146 -415
rect -112 -449 -106 -415
rect -152 -487 -106 -449
rect -152 -521 -146 -487
rect -112 -521 -106 -487
rect -152 -536 -106 -521
rect 106 449 152 464
rect 106 415 112 449
rect 146 415 152 449
rect 106 377 152 415
rect 106 343 112 377
rect 146 343 152 377
rect 106 305 152 343
rect 106 271 112 305
rect 146 271 152 305
rect 106 233 152 271
rect 106 199 112 233
rect 146 199 152 233
rect 106 161 152 199
rect 106 127 112 161
rect 146 127 152 161
rect 106 89 152 127
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -127 152 -89
rect 106 -161 112 -127
rect 146 -161 152 -127
rect 106 -199 152 -161
rect 106 -233 112 -199
rect 146 -233 152 -199
rect 106 -271 152 -233
rect 106 -305 112 -271
rect 146 -305 152 -271
rect 106 -343 152 -305
rect 106 -377 112 -343
rect 146 -377 152 -343
rect 106 -415 152 -377
rect 106 -449 112 -415
rect 146 -449 152 -415
rect 106 -487 152 -449
rect 106 -521 112 -487
rect 146 -521 152 -487
rect 106 -536 152 -521
<< end >>
