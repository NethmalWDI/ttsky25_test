magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -823 4997 6783 5083
rect -823 -587 -737 4997
rect 1794 4776 1946 4806
rect 1794 4664 1966 4776
rect 6697 -587 6783 4997
rect -823 -673 6783 -587
<< nmoslvt >>
rect 1820 4750 1920 4780
rect 1820 4690 1940 4750
<< psubdiff >>
rect -797 5023 -709 5057
rect -675 5023 -641 5057
rect -607 5023 -573 5057
rect -539 5023 -505 5057
rect -471 5023 -437 5057
rect -403 5023 -369 5057
rect -335 5023 -301 5057
rect -267 5023 -233 5057
rect -199 5023 -165 5057
rect -131 5023 -97 5057
rect -63 5023 -29 5057
rect 5 5023 39 5057
rect 73 5023 107 5057
rect 141 5023 175 5057
rect 209 5023 243 5057
rect 277 5023 311 5057
rect 345 5023 379 5057
rect 413 5023 447 5057
rect 481 5023 515 5057
rect 549 5023 583 5057
rect 617 5023 651 5057
rect 685 5023 719 5057
rect 753 5023 787 5057
rect 821 5023 855 5057
rect 889 5023 923 5057
rect 957 5023 991 5057
rect 1025 5023 1059 5057
rect 1093 5023 1127 5057
rect 1161 5023 1195 5057
rect 1229 5023 1263 5057
rect 1297 5023 1331 5057
rect 1365 5023 1399 5057
rect 1433 5023 1467 5057
rect 1501 5023 1535 5057
rect 1569 5023 1603 5057
rect 1637 5023 1671 5057
rect 1705 5023 1739 5057
rect 1773 5023 1807 5057
rect 1841 5023 1875 5057
rect 1909 5023 1943 5057
rect 1977 5023 2011 5057
rect 2045 5023 2079 5057
rect 2113 5023 2147 5057
rect 2181 5023 2215 5057
rect 2249 5023 2283 5057
rect 2317 5023 2351 5057
rect 2385 5023 2419 5057
rect 2453 5023 2487 5057
rect 2521 5023 2555 5057
rect 2589 5023 2623 5057
rect 2657 5023 2691 5057
rect 2725 5023 2759 5057
rect 2793 5023 2827 5057
rect 2861 5023 2895 5057
rect 2929 5023 2963 5057
rect 2997 5023 3031 5057
rect 3065 5023 3099 5057
rect 3133 5023 3167 5057
rect 3201 5023 3235 5057
rect 3269 5023 3303 5057
rect 3337 5023 3371 5057
rect 3405 5023 3439 5057
rect 3473 5023 3507 5057
rect 3541 5023 3575 5057
rect 3609 5023 3643 5057
rect 3677 5023 3711 5057
rect 3745 5023 3779 5057
rect 3813 5023 3847 5057
rect 3881 5023 3915 5057
rect 3949 5023 3983 5057
rect 4017 5023 4051 5057
rect 4085 5023 4119 5057
rect 4153 5023 4187 5057
rect 4221 5023 4255 5057
rect 4289 5023 4323 5057
rect 4357 5023 4391 5057
rect 4425 5023 4459 5057
rect 4493 5023 4527 5057
rect 4561 5023 4595 5057
rect 4629 5023 4663 5057
rect 4697 5023 4731 5057
rect 4765 5023 4799 5057
rect 4833 5023 4867 5057
rect 4901 5023 4935 5057
rect 4969 5023 5003 5057
rect 5037 5023 5071 5057
rect 5105 5023 5139 5057
rect 5173 5023 5207 5057
rect 5241 5023 5275 5057
rect 5309 5023 5343 5057
rect 5377 5023 5411 5057
rect 5445 5023 5479 5057
rect 5513 5023 5547 5057
rect 5581 5023 5615 5057
rect 5649 5023 5683 5057
rect 5717 5023 5751 5057
rect 5785 5023 5819 5057
rect 5853 5023 5887 5057
rect 5921 5023 5955 5057
rect 5989 5023 6023 5057
rect 6057 5023 6091 5057
rect 6125 5023 6159 5057
rect 6193 5023 6227 5057
rect 6261 5023 6295 5057
rect 6329 5023 6363 5057
rect 6397 5023 6431 5057
rect 6465 5023 6499 5057
rect 6533 5023 6567 5057
rect 6601 5023 6635 5057
rect 6669 5023 6757 5057
rect -797 4976 -763 5023
rect -797 4908 -763 4942
rect -797 4840 -763 4874
rect -797 4772 -763 4806
rect 6723 4976 6757 5023
rect 6723 4908 6757 4942
rect 6723 4840 6757 4874
rect -797 4704 -763 4738
rect 6723 4772 6757 4806
rect 6723 4704 6757 4738
rect -797 4636 -763 4670
rect -797 4568 -763 4602
rect -797 4500 -763 4534
rect -797 4432 -763 4466
rect -797 4364 -763 4398
rect -797 4296 -763 4330
rect -797 4228 -763 4262
rect -797 4160 -763 4194
rect -797 4092 -763 4126
rect -797 4024 -763 4058
rect -797 3956 -763 3990
rect -797 3888 -763 3922
rect -797 3820 -763 3854
rect -797 3752 -763 3786
rect -797 3684 -763 3718
rect -797 3616 -763 3650
rect -797 3548 -763 3582
rect -797 3480 -763 3514
rect -797 3412 -763 3446
rect -797 3344 -763 3378
rect -797 3276 -763 3310
rect -797 3208 -763 3242
rect -797 3140 -763 3174
rect -797 3072 -763 3106
rect -797 3004 -763 3038
rect -797 2936 -763 2970
rect -797 2868 -763 2902
rect -797 2800 -763 2834
rect -797 2732 -763 2766
rect -797 2664 -763 2698
rect -797 2596 -763 2630
rect -797 2528 -763 2562
rect -797 2460 -763 2494
rect -797 2392 -763 2426
rect -797 2324 -763 2358
rect -797 2256 -763 2290
rect -797 2188 -763 2222
rect -797 2120 -763 2154
rect -797 2052 -763 2086
rect -797 1984 -763 2018
rect -797 1916 -763 1950
rect -797 1848 -763 1882
rect -797 1780 -763 1814
rect -797 1712 -763 1746
rect -797 1644 -763 1678
rect -797 1576 -763 1610
rect -797 1508 -763 1542
rect -797 1440 -763 1474
rect -797 1372 -763 1406
rect -797 1304 -763 1338
rect -797 1236 -763 1270
rect -797 1168 -763 1202
rect -797 1100 -763 1134
rect -797 1032 -763 1066
rect -797 964 -763 998
rect -797 896 -763 930
rect -797 828 -763 862
rect -797 760 -763 794
rect -797 692 -763 726
rect -797 624 -763 658
rect -797 556 -763 590
rect -797 488 -763 522
rect -797 420 -763 454
rect -797 352 -763 386
rect -797 284 -763 318
rect -797 216 -763 250
rect -797 148 -763 182
rect -797 80 -763 114
rect -797 12 -763 46
rect -797 -56 -763 -22
rect -797 -124 -763 -90
rect -797 -192 -763 -158
rect -797 -260 -763 -226
rect -797 -328 -763 -294
rect -797 -396 -763 -362
rect -797 -464 -763 -430
rect -797 -532 -763 -498
rect -797 -613 -763 -566
rect 6723 4636 6757 4670
rect 6723 4568 6757 4602
rect 6723 4500 6757 4534
rect 6723 4432 6757 4466
rect 6723 4364 6757 4398
rect 6723 4296 6757 4330
rect 6723 4228 6757 4262
rect 6723 4160 6757 4194
rect 6723 4092 6757 4126
rect 6723 4024 6757 4058
rect 6723 3956 6757 3990
rect 6723 3888 6757 3922
rect 6723 3820 6757 3854
rect 6723 3752 6757 3786
rect 6723 3684 6757 3718
rect 6723 3616 6757 3650
rect 6723 3548 6757 3582
rect 6723 3480 6757 3514
rect 6723 3412 6757 3446
rect 6723 3344 6757 3378
rect 6723 3276 6757 3310
rect 6723 3208 6757 3242
rect 6723 3140 6757 3174
rect 6723 3072 6757 3106
rect 6723 3004 6757 3038
rect 6723 2936 6757 2970
rect 6723 2868 6757 2902
rect 6723 2800 6757 2834
rect 6723 2732 6757 2766
rect 6723 2664 6757 2698
rect 6723 2596 6757 2630
rect 6723 2528 6757 2562
rect 6723 2460 6757 2494
rect 6723 2392 6757 2426
rect 6723 2324 6757 2358
rect 6723 2256 6757 2290
rect 6723 2188 6757 2222
rect 6723 2120 6757 2154
rect 6723 2052 6757 2086
rect 6723 1984 6757 2018
rect 6723 1916 6757 1950
rect 6723 1848 6757 1882
rect 6723 1780 6757 1814
rect 6723 1712 6757 1746
rect 6723 1644 6757 1678
rect 6723 1576 6757 1610
rect 6723 1508 6757 1542
rect 6723 1440 6757 1474
rect 6723 1372 6757 1406
rect 6723 1304 6757 1338
rect 6723 1236 6757 1270
rect 6723 1168 6757 1202
rect 6723 1100 6757 1134
rect 6723 1032 6757 1066
rect 6723 964 6757 998
rect 6723 896 6757 930
rect 6723 828 6757 862
rect 6723 760 6757 794
rect 6723 692 6757 726
rect 6723 624 6757 658
rect 6723 556 6757 590
rect 6723 488 6757 522
rect 6723 420 6757 454
rect 6723 352 6757 386
rect 6723 284 6757 318
rect 6723 216 6757 250
rect 6723 148 6757 182
rect 6723 80 6757 114
rect 6723 12 6757 46
rect 6723 -56 6757 -22
rect 6723 -124 6757 -90
rect 6723 -192 6757 -158
rect 6723 -260 6757 -226
rect 6723 -328 6757 -294
rect 6723 -396 6757 -362
rect 6723 -464 6757 -430
rect 6723 -532 6757 -498
rect 6723 -613 6757 -566
rect -797 -647 -709 -613
rect -675 -647 -641 -613
rect -607 -647 -573 -613
rect -539 -647 -505 -613
rect -471 -647 -437 -613
rect -403 -647 -369 -613
rect -335 -647 -301 -613
rect -267 -647 -233 -613
rect -199 -647 -165 -613
rect -131 -647 -97 -613
rect -63 -647 -29 -613
rect 5 -647 39 -613
rect 73 -647 107 -613
rect 141 -647 175 -613
rect 209 -647 243 -613
rect 277 -647 311 -613
rect 345 -647 379 -613
rect 413 -647 447 -613
rect 481 -647 515 -613
rect 549 -647 583 -613
rect 617 -647 651 -613
rect 685 -647 719 -613
rect 753 -647 787 -613
rect 821 -647 855 -613
rect 889 -647 923 -613
rect 957 -647 991 -613
rect 1025 -647 1059 -613
rect 1093 -647 1127 -613
rect 1161 -647 1195 -613
rect 1229 -647 1263 -613
rect 1297 -647 1331 -613
rect 1365 -647 1399 -613
rect 1433 -647 1467 -613
rect 1501 -647 1535 -613
rect 1569 -647 1603 -613
rect 1637 -647 1671 -613
rect 1705 -647 1739 -613
rect 1773 -647 1807 -613
rect 1841 -647 1875 -613
rect 1909 -647 1943 -613
rect 1977 -647 2011 -613
rect 2045 -647 2079 -613
rect 2113 -647 2147 -613
rect 2181 -647 2215 -613
rect 2249 -647 2283 -613
rect 2317 -647 2351 -613
rect 2385 -647 2419 -613
rect 2453 -647 2487 -613
rect 2521 -647 2555 -613
rect 2589 -647 2623 -613
rect 2657 -647 2691 -613
rect 2725 -647 2759 -613
rect 2793 -647 2827 -613
rect 2861 -647 2895 -613
rect 2929 -647 2963 -613
rect 2997 -647 3031 -613
rect 3065 -647 3099 -613
rect 3133 -647 3167 -613
rect 3201 -647 3235 -613
rect 3269 -647 3303 -613
rect 3337 -647 3371 -613
rect 3405 -647 3439 -613
rect 3473 -647 3507 -613
rect 3541 -647 3575 -613
rect 3609 -647 3643 -613
rect 3677 -647 3711 -613
rect 3745 -647 3779 -613
rect 3813 -647 3847 -613
rect 3881 -647 3915 -613
rect 3949 -647 3983 -613
rect 4017 -647 4051 -613
rect 4085 -647 4119 -613
rect 4153 -647 4187 -613
rect 4221 -647 4255 -613
rect 4289 -647 4323 -613
rect 4357 -647 4391 -613
rect 4425 -647 4459 -613
rect 4493 -647 4527 -613
rect 4561 -647 4595 -613
rect 4629 -647 4663 -613
rect 4697 -647 4731 -613
rect 4765 -647 4799 -613
rect 4833 -647 4867 -613
rect 4901 -647 4935 -613
rect 4969 -647 5003 -613
rect 5037 -647 5071 -613
rect 5105 -647 5139 -613
rect 5173 -647 5207 -613
rect 5241 -647 5275 -613
rect 5309 -647 5343 -613
rect 5377 -647 5411 -613
rect 5445 -647 5479 -613
rect 5513 -647 5547 -613
rect 5581 -647 5615 -613
rect 5649 -647 5683 -613
rect 5717 -647 5751 -613
rect 5785 -647 5819 -613
rect 5853 -647 5887 -613
rect 5921 -647 5955 -613
rect 5989 -647 6023 -613
rect 6057 -647 6091 -613
rect 6125 -647 6159 -613
rect 6193 -647 6227 -613
rect 6261 -647 6295 -613
rect 6329 -647 6363 -613
rect 6397 -647 6431 -613
rect 6465 -647 6499 -613
rect 6533 -647 6567 -613
rect 6601 -647 6635 -613
rect 6669 -647 6757 -613
<< psubdiffcont >>
rect -709 5023 -675 5057
rect -641 5023 -607 5057
rect -573 5023 -539 5057
rect -505 5023 -471 5057
rect -437 5023 -403 5057
rect -369 5023 -335 5057
rect -301 5023 -267 5057
rect -233 5023 -199 5057
rect -165 5023 -131 5057
rect -97 5023 -63 5057
rect -29 5023 5 5057
rect 39 5023 73 5057
rect 107 5023 141 5057
rect 175 5023 209 5057
rect 243 5023 277 5057
rect 311 5023 345 5057
rect 379 5023 413 5057
rect 447 5023 481 5057
rect 515 5023 549 5057
rect 583 5023 617 5057
rect 651 5023 685 5057
rect 719 5023 753 5057
rect 787 5023 821 5057
rect 855 5023 889 5057
rect 923 5023 957 5057
rect 991 5023 1025 5057
rect 1059 5023 1093 5057
rect 1127 5023 1161 5057
rect 1195 5023 1229 5057
rect 1263 5023 1297 5057
rect 1331 5023 1365 5057
rect 1399 5023 1433 5057
rect 1467 5023 1501 5057
rect 1535 5023 1569 5057
rect 1603 5023 1637 5057
rect 1671 5023 1705 5057
rect 1739 5023 1773 5057
rect 1807 5023 1841 5057
rect 1875 5023 1909 5057
rect 1943 5023 1977 5057
rect 2011 5023 2045 5057
rect 2079 5023 2113 5057
rect 2147 5023 2181 5057
rect 2215 5023 2249 5057
rect 2283 5023 2317 5057
rect 2351 5023 2385 5057
rect 2419 5023 2453 5057
rect 2487 5023 2521 5057
rect 2555 5023 2589 5057
rect 2623 5023 2657 5057
rect 2691 5023 2725 5057
rect 2759 5023 2793 5057
rect 2827 5023 2861 5057
rect 2895 5023 2929 5057
rect 2963 5023 2997 5057
rect 3031 5023 3065 5057
rect 3099 5023 3133 5057
rect 3167 5023 3201 5057
rect 3235 5023 3269 5057
rect 3303 5023 3337 5057
rect 3371 5023 3405 5057
rect 3439 5023 3473 5057
rect 3507 5023 3541 5057
rect 3575 5023 3609 5057
rect 3643 5023 3677 5057
rect 3711 5023 3745 5057
rect 3779 5023 3813 5057
rect 3847 5023 3881 5057
rect 3915 5023 3949 5057
rect 3983 5023 4017 5057
rect 4051 5023 4085 5057
rect 4119 5023 4153 5057
rect 4187 5023 4221 5057
rect 4255 5023 4289 5057
rect 4323 5023 4357 5057
rect 4391 5023 4425 5057
rect 4459 5023 4493 5057
rect 4527 5023 4561 5057
rect 4595 5023 4629 5057
rect 4663 5023 4697 5057
rect 4731 5023 4765 5057
rect 4799 5023 4833 5057
rect 4867 5023 4901 5057
rect 4935 5023 4969 5057
rect 5003 5023 5037 5057
rect 5071 5023 5105 5057
rect 5139 5023 5173 5057
rect 5207 5023 5241 5057
rect 5275 5023 5309 5057
rect 5343 5023 5377 5057
rect 5411 5023 5445 5057
rect 5479 5023 5513 5057
rect 5547 5023 5581 5057
rect 5615 5023 5649 5057
rect 5683 5023 5717 5057
rect 5751 5023 5785 5057
rect 5819 5023 5853 5057
rect 5887 5023 5921 5057
rect 5955 5023 5989 5057
rect 6023 5023 6057 5057
rect 6091 5023 6125 5057
rect 6159 5023 6193 5057
rect 6227 5023 6261 5057
rect 6295 5023 6329 5057
rect 6363 5023 6397 5057
rect 6431 5023 6465 5057
rect 6499 5023 6533 5057
rect 6567 5023 6601 5057
rect 6635 5023 6669 5057
rect -797 4942 -763 4976
rect -797 4874 -763 4908
rect -797 4806 -763 4840
rect 6723 4942 6757 4976
rect 6723 4874 6757 4908
rect 6723 4806 6757 4840
rect -797 4738 -763 4772
rect -797 4670 -763 4704
rect 6723 4738 6757 4772
rect -797 4602 -763 4636
rect -797 4534 -763 4568
rect -797 4466 -763 4500
rect -797 4398 -763 4432
rect -797 4330 -763 4364
rect -797 4262 -763 4296
rect -797 4194 -763 4228
rect -797 4126 -763 4160
rect -797 4058 -763 4092
rect -797 3990 -763 4024
rect -797 3922 -763 3956
rect -797 3854 -763 3888
rect -797 3786 -763 3820
rect -797 3718 -763 3752
rect -797 3650 -763 3684
rect -797 3582 -763 3616
rect -797 3514 -763 3548
rect -797 3446 -763 3480
rect -797 3378 -763 3412
rect -797 3310 -763 3344
rect -797 3242 -763 3276
rect -797 3174 -763 3208
rect -797 3106 -763 3140
rect -797 3038 -763 3072
rect -797 2970 -763 3004
rect -797 2902 -763 2936
rect -797 2834 -763 2868
rect -797 2766 -763 2800
rect -797 2698 -763 2732
rect -797 2630 -763 2664
rect -797 2562 -763 2596
rect -797 2494 -763 2528
rect -797 2426 -763 2460
rect -797 2358 -763 2392
rect -797 2290 -763 2324
rect -797 2222 -763 2256
rect -797 2154 -763 2188
rect -797 2086 -763 2120
rect -797 2018 -763 2052
rect -797 1950 -763 1984
rect -797 1882 -763 1916
rect -797 1814 -763 1848
rect -797 1746 -763 1780
rect -797 1678 -763 1712
rect -797 1610 -763 1644
rect -797 1542 -763 1576
rect -797 1474 -763 1508
rect -797 1406 -763 1440
rect -797 1338 -763 1372
rect -797 1270 -763 1304
rect -797 1202 -763 1236
rect -797 1134 -763 1168
rect -797 1066 -763 1100
rect -797 998 -763 1032
rect -797 930 -763 964
rect -797 862 -763 896
rect -797 794 -763 828
rect -797 726 -763 760
rect -797 658 -763 692
rect -797 590 -763 624
rect -797 522 -763 556
rect -797 454 -763 488
rect -797 386 -763 420
rect -797 318 -763 352
rect -797 250 -763 284
rect -797 182 -763 216
rect -797 114 -763 148
rect -797 46 -763 80
rect -797 -22 -763 12
rect -797 -90 -763 -56
rect -797 -158 -763 -124
rect -797 -226 -763 -192
rect -797 -294 -763 -260
rect -797 -362 -763 -328
rect -797 -430 -763 -396
rect -797 -498 -763 -464
rect -797 -566 -763 -532
rect 6723 4670 6757 4704
rect 6723 4602 6757 4636
rect 6723 4534 6757 4568
rect 6723 4466 6757 4500
rect 6723 4398 6757 4432
rect 6723 4330 6757 4364
rect 6723 4262 6757 4296
rect 6723 4194 6757 4228
rect 6723 4126 6757 4160
rect 6723 4058 6757 4092
rect 6723 3990 6757 4024
rect 6723 3922 6757 3956
rect 6723 3854 6757 3888
rect 6723 3786 6757 3820
rect 6723 3718 6757 3752
rect 6723 3650 6757 3684
rect 6723 3582 6757 3616
rect 6723 3514 6757 3548
rect 6723 3446 6757 3480
rect 6723 3378 6757 3412
rect 6723 3310 6757 3344
rect 6723 3242 6757 3276
rect 6723 3174 6757 3208
rect 6723 3106 6757 3140
rect 6723 3038 6757 3072
rect 6723 2970 6757 3004
rect 6723 2902 6757 2936
rect 6723 2834 6757 2868
rect 6723 2766 6757 2800
rect 6723 2698 6757 2732
rect 6723 2630 6757 2664
rect 6723 2562 6757 2596
rect 6723 2494 6757 2528
rect 6723 2426 6757 2460
rect 6723 2358 6757 2392
rect 6723 2290 6757 2324
rect 6723 2222 6757 2256
rect 6723 2154 6757 2188
rect 6723 2086 6757 2120
rect 6723 2018 6757 2052
rect 6723 1950 6757 1984
rect 6723 1882 6757 1916
rect 6723 1814 6757 1848
rect 6723 1746 6757 1780
rect 6723 1678 6757 1712
rect 6723 1610 6757 1644
rect 6723 1542 6757 1576
rect 6723 1474 6757 1508
rect 6723 1406 6757 1440
rect 6723 1338 6757 1372
rect 6723 1270 6757 1304
rect 6723 1202 6757 1236
rect 6723 1134 6757 1168
rect 6723 1066 6757 1100
rect 6723 998 6757 1032
rect 6723 930 6757 964
rect 6723 862 6757 896
rect 6723 794 6757 828
rect 6723 726 6757 760
rect 6723 658 6757 692
rect 6723 590 6757 624
rect 6723 522 6757 556
rect 6723 454 6757 488
rect 6723 386 6757 420
rect 6723 318 6757 352
rect 6723 250 6757 284
rect 6723 182 6757 216
rect 6723 114 6757 148
rect 6723 46 6757 80
rect 6723 -22 6757 12
rect 6723 -90 6757 -56
rect 6723 -158 6757 -124
rect 6723 -226 6757 -192
rect 6723 -294 6757 -260
rect 6723 -362 6757 -328
rect 6723 -430 6757 -396
rect 6723 -498 6757 -464
rect 6723 -566 6757 -532
rect -709 -647 -675 -613
rect -641 -647 -607 -613
rect -573 -647 -539 -613
rect -505 -647 -471 -613
rect -437 -647 -403 -613
rect -369 -647 -335 -613
rect -301 -647 -267 -613
rect -233 -647 -199 -613
rect -165 -647 -131 -613
rect -97 -647 -63 -613
rect -29 -647 5 -613
rect 39 -647 73 -613
rect 107 -647 141 -613
rect 175 -647 209 -613
rect 243 -647 277 -613
rect 311 -647 345 -613
rect 379 -647 413 -613
rect 447 -647 481 -613
rect 515 -647 549 -613
rect 583 -647 617 -613
rect 651 -647 685 -613
rect 719 -647 753 -613
rect 787 -647 821 -613
rect 855 -647 889 -613
rect 923 -647 957 -613
rect 991 -647 1025 -613
rect 1059 -647 1093 -613
rect 1127 -647 1161 -613
rect 1195 -647 1229 -613
rect 1263 -647 1297 -613
rect 1331 -647 1365 -613
rect 1399 -647 1433 -613
rect 1467 -647 1501 -613
rect 1535 -647 1569 -613
rect 1603 -647 1637 -613
rect 1671 -647 1705 -613
rect 1739 -647 1773 -613
rect 1807 -647 1841 -613
rect 1875 -647 1909 -613
rect 1943 -647 1977 -613
rect 2011 -647 2045 -613
rect 2079 -647 2113 -613
rect 2147 -647 2181 -613
rect 2215 -647 2249 -613
rect 2283 -647 2317 -613
rect 2351 -647 2385 -613
rect 2419 -647 2453 -613
rect 2487 -647 2521 -613
rect 2555 -647 2589 -613
rect 2623 -647 2657 -613
rect 2691 -647 2725 -613
rect 2759 -647 2793 -613
rect 2827 -647 2861 -613
rect 2895 -647 2929 -613
rect 2963 -647 2997 -613
rect 3031 -647 3065 -613
rect 3099 -647 3133 -613
rect 3167 -647 3201 -613
rect 3235 -647 3269 -613
rect 3303 -647 3337 -613
rect 3371 -647 3405 -613
rect 3439 -647 3473 -613
rect 3507 -647 3541 -613
rect 3575 -647 3609 -613
rect 3643 -647 3677 -613
rect 3711 -647 3745 -613
rect 3779 -647 3813 -613
rect 3847 -647 3881 -613
rect 3915 -647 3949 -613
rect 3983 -647 4017 -613
rect 4051 -647 4085 -613
rect 4119 -647 4153 -613
rect 4187 -647 4221 -613
rect 4255 -647 4289 -613
rect 4323 -647 4357 -613
rect 4391 -647 4425 -613
rect 4459 -647 4493 -613
rect 4527 -647 4561 -613
rect 4595 -647 4629 -613
rect 4663 -647 4697 -613
rect 4731 -647 4765 -613
rect 4799 -647 4833 -613
rect 4867 -647 4901 -613
rect 4935 -647 4969 -613
rect 5003 -647 5037 -613
rect 5071 -647 5105 -613
rect 5139 -647 5173 -613
rect 5207 -647 5241 -613
rect 5275 -647 5309 -613
rect 5343 -647 5377 -613
rect 5411 -647 5445 -613
rect 5479 -647 5513 -613
rect 5547 -647 5581 -613
rect 5615 -647 5649 -613
rect 5683 -647 5717 -613
rect 5751 -647 5785 -613
rect 5819 -647 5853 -613
rect 5887 -647 5921 -613
rect 5955 -647 5989 -613
rect 6023 -647 6057 -613
rect 6091 -647 6125 -613
rect 6159 -647 6193 -613
rect 6227 -647 6261 -613
rect 6295 -647 6329 -613
rect 6363 -647 6397 -613
rect 6431 -647 6465 -613
rect 6499 -647 6533 -613
rect 6567 -647 6601 -613
rect 6635 -647 6669 -613
<< locali >>
rect -797 5023 -709 5057
rect -675 5023 -641 5057
rect -607 5023 -573 5057
rect -539 5023 -505 5057
rect -471 5023 -437 5057
rect -403 5023 -369 5057
rect -335 5023 -301 5057
rect -267 5023 -233 5057
rect -199 5023 -165 5057
rect -131 5023 -97 5057
rect -63 5023 -29 5057
rect 5 5023 39 5057
rect 73 5023 107 5057
rect 141 5023 175 5057
rect 209 5023 243 5057
rect 277 5023 311 5057
rect 345 5023 379 5057
rect 413 5023 447 5057
rect 481 5023 515 5057
rect 549 5023 583 5057
rect 617 5023 651 5057
rect 685 5023 719 5057
rect 753 5023 787 5057
rect 821 5023 855 5057
rect 889 5023 923 5057
rect 957 5023 991 5057
rect 1025 5023 1059 5057
rect 1093 5023 1127 5057
rect 1161 5023 1195 5057
rect 1229 5023 1263 5057
rect 1297 5023 1331 5057
rect 1365 5023 1399 5057
rect 1433 5023 1467 5057
rect 1501 5023 1535 5057
rect 1569 5023 1603 5057
rect 1637 5023 1671 5057
rect 1705 5023 1739 5057
rect 1773 5023 1807 5057
rect 1841 5023 1875 5057
rect 1909 5023 1943 5057
rect 1977 5023 2011 5057
rect 2045 5023 2079 5057
rect 2113 5023 2147 5057
rect 2181 5023 2215 5057
rect 2249 5023 2283 5057
rect 2317 5023 2351 5057
rect 2385 5023 2419 5057
rect 2453 5023 2487 5057
rect 2521 5023 2555 5057
rect 2589 5023 2623 5057
rect 2657 5023 2691 5057
rect 2725 5023 2759 5057
rect 2793 5023 2827 5057
rect 2861 5023 2895 5057
rect 2929 5023 2963 5057
rect 2997 5023 3031 5057
rect 3065 5023 3099 5057
rect 3133 5023 3167 5057
rect 3201 5023 3235 5057
rect 3269 5023 3303 5057
rect 3337 5023 3371 5057
rect 3405 5023 3439 5057
rect 3473 5023 3507 5057
rect 3541 5023 3575 5057
rect 3609 5023 3643 5057
rect 3677 5023 3711 5057
rect 3745 5023 3779 5057
rect 3813 5023 3847 5057
rect 3881 5023 3915 5057
rect 3949 5023 3983 5057
rect 4017 5023 4051 5057
rect 4085 5023 4119 5057
rect 4153 5023 4187 5057
rect 4221 5023 4255 5057
rect 4289 5023 4323 5057
rect 4357 5023 4391 5057
rect 4425 5023 4459 5057
rect 4493 5023 4527 5057
rect 4561 5023 4595 5057
rect 4629 5023 4663 5057
rect 4697 5023 4731 5057
rect 4765 5023 4799 5057
rect 4833 5023 4867 5057
rect 4901 5023 4935 5057
rect 4969 5023 5003 5057
rect 5037 5023 5071 5057
rect 5105 5023 5139 5057
rect 5173 5023 5207 5057
rect 5241 5023 5275 5057
rect 5309 5023 5343 5057
rect 5377 5023 5411 5057
rect 5445 5023 5479 5057
rect 5513 5023 5547 5057
rect 5581 5023 5615 5057
rect 5649 5023 5683 5057
rect 5717 5023 5751 5057
rect 5785 5023 5819 5057
rect 5853 5023 5887 5057
rect 5921 5023 5955 5057
rect 5989 5023 6023 5057
rect 6057 5023 6091 5057
rect 6125 5023 6159 5057
rect 6193 5023 6227 5057
rect 6261 5023 6295 5057
rect 6329 5023 6363 5057
rect 6397 5023 6431 5057
rect 6465 5023 6499 5057
rect 6533 5023 6567 5057
rect 6601 5023 6635 5057
rect 6669 5023 6757 5057
rect -797 4976 -763 5023
rect -797 4908 -763 4942
rect -797 4840 -763 4874
rect -797 4772 -763 4806
rect -797 4704 -763 4738
rect -797 4636 -763 4670
rect -797 4568 -763 4602
rect -797 4500 -763 4534
rect -797 4432 -763 4466
rect -797 4364 -763 4398
rect -797 4296 -763 4330
rect -797 4228 -763 4262
rect -797 4160 -763 4194
rect -797 4092 -763 4126
rect -797 4024 -763 4058
rect -797 3956 -763 3990
rect -797 3888 -763 3922
rect -797 3820 -763 3854
rect -797 3752 -763 3786
rect -797 3684 -763 3718
rect -797 3616 -763 3650
rect -797 3548 -763 3582
rect -797 3480 -763 3514
rect -797 3412 -763 3446
rect -797 3344 -763 3378
rect -797 3276 -763 3310
rect -797 3208 -763 3242
rect -797 3140 -763 3174
rect -797 3072 -763 3106
rect -797 3004 -763 3038
rect -797 2936 -763 2970
rect -797 2868 -763 2902
rect -797 2800 -763 2834
rect -797 2732 -763 2766
rect -797 2664 -763 2698
rect -797 2596 -763 2630
rect -797 2528 -763 2562
rect -797 2460 -763 2494
rect -797 2392 -763 2426
rect -797 2324 -763 2358
rect -797 2256 -763 2290
rect -797 2188 -763 2222
rect -797 2120 -763 2154
rect -797 2052 -763 2086
rect -797 1984 -763 2018
rect -797 1916 -763 1950
rect -797 1848 -763 1882
rect -797 1780 -763 1814
rect -797 1712 -763 1746
rect -797 1644 -763 1678
rect -797 1576 -763 1610
rect -797 1508 -763 1542
rect -797 1440 -763 1474
rect -797 1372 -763 1406
rect -797 1304 -763 1338
rect -797 1236 -763 1270
rect -797 1168 -763 1202
rect -797 1100 -763 1134
rect -797 1032 -763 1066
rect -797 964 -763 998
rect -797 896 -763 930
rect -797 828 -763 862
rect -797 760 -763 794
rect -797 692 -763 726
rect -797 624 -763 658
rect -797 556 -763 590
rect -797 488 -763 522
rect -797 420 -763 454
rect -797 352 -763 386
rect -797 284 -763 318
rect -797 216 -763 250
rect -797 148 -763 182
rect -797 80 -763 114
rect -797 12 -763 46
rect -797 -56 -763 -22
rect -797 -124 -763 -90
rect -797 -192 -763 -158
rect -797 -260 -763 -226
rect -797 -328 -763 -294
rect -797 -396 -763 -362
rect -797 -464 -763 -430
rect -797 -532 -763 -498
rect -797 -613 -763 -566
rect 6723 4976 6757 5023
rect 6723 4908 6757 4942
rect 6723 4840 6757 4874
rect 6723 4772 6757 4806
rect 6723 4704 6757 4738
rect 6723 4636 6757 4670
rect 6723 4568 6757 4602
rect 6723 4500 6757 4534
rect 6723 4432 6757 4466
rect 6723 4364 6757 4398
rect 6723 4296 6757 4330
rect 6723 4228 6757 4262
rect 6723 4160 6757 4194
rect 6723 4092 6757 4126
rect 6723 4024 6757 4058
rect 6723 3956 6757 3990
rect 6723 3888 6757 3922
rect 6723 3820 6757 3854
rect 6723 3752 6757 3786
rect 6723 3684 6757 3718
rect 6723 3616 6757 3650
rect 6723 3548 6757 3582
rect 6723 3480 6757 3514
rect 6723 3412 6757 3446
rect 6723 3344 6757 3378
rect 6723 3276 6757 3310
rect 6723 3208 6757 3242
rect 6723 3140 6757 3174
rect 6723 3072 6757 3106
rect 6723 3004 6757 3038
rect 6723 2936 6757 2970
rect 6723 2868 6757 2902
rect 6723 2800 6757 2834
rect 6723 2732 6757 2766
rect 6723 2664 6757 2698
rect 6723 2596 6757 2630
rect 6723 2528 6757 2562
rect 6723 2460 6757 2494
rect 6723 2392 6757 2426
rect 6723 2324 6757 2358
rect 6723 2256 6757 2290
rect 6723 2188 6757 2222
rect 6723 2120 6757 2154
rect 6723 2052 6757 2086
rect 6723 1984 6757 2018
rect 6723 1916 6757 1950
rect 6723 1848 6757 1882
rect 6723 1780 6757 1814
rect 6723 1712 6757 1746
rect 6723 1644 6757 1678
rect 6723 1576 6757 1610
rect 6723 1508 6757 1542
rect 6723 1440 6757 1474
rect 6723 1372 6757 1406
rect 6723 1304 6757 1338
rect 6723 1236 6757 1270
rect 6723 1168 6757 1202
rect 6723 1100 6757 1134
rect 6723 1032 6757 1066
rect 6723 964 6757 998
rect 6723 896 6757 930
rect 6723 828 6757 862
rect 6723 760 6757 794
rect 6723 692 6757 726
rect 6723 624 6757 658
rect 6723 556 6757 590
rect 6723 488 6757 522
rect 6723 420 6757 454
rect 6723 352 6757 386
rect 6723 284 6757 318
rect 6723 216 6757 250
rect 6723 148 6757 182
rect 6723 80 6757 114
rect 6723 12 6757 46
rect 6723 -56 6757 -22
rect 6723 -124 6757 -90
rect 6723 -192 6757 -158
rect 6723 -260 6757 -226
rect 6723 -328 6757 -294
rect 6723 -396 6757 -362
rect 6723 -464 6757 -430
rect 6723 -532 6757 -498
rect 6723 -613 6757 -566
rect -797 -647 -709 -613
rect -675 -647 -641 -613
rect -607 -647 -573 -613
rect -539 -647 -505 -613
rect -471 -647 -437 -613
rect -403 -647 -369 -613
rect -335 -647 -301 -613
rect -267 -647 -233 -613
rect -199 -647 -165 -613
rect -131 -647 -97 -613
rect -63 -647 -29 -613
rect 5 -647 39 -613
rect 73 -647 107 -613
rect 141 -647 175 -613
rect 209 -647 243 -613
rect 277 -647 311 -613
rect 345 -647 379 -613
rect 413 -647 447 -613
rect 481 -647 515 -613
rect 549 -647 583 -613
rect 617 -647 651 -613
rect 685 -647 719 -613
rect 753 -647 787 -613
rect 821 -647 855 -613
rect 889 -647 923 -613
rect 957 -647 991 -613
rect 1025 -647 1059 -613
rect 1093 -647 1127 -613
rect 1161 -647 1195 -613
rect 1229 -647 1263 -613
rect 1297 -647 1331 -613
rect 1365 -647 1399 -613
rect 1433 -647 1467 -613
rect 1501 -647 1535 -613
rect 1569 -647 1603 -613
rect 1637 -647 1671 -613
rect 1705 -647 1739 -613
rect 1773 -647 1807 -613
rect 1841 -647 1875 -613
rect 1909 -647 1943 -613
rect 1977 -647 2011 -613
rect 2045 -647 2079 -613
rect 2113 -647 2147 -613
rect 2181 -647 2215 -613
rect 2249 -647 2283 -613
rect 2317 -647 2351 -613
rect 2385 -647 2419 -613
rect 2453 -647 2487 -613
rect 2521 -647 2555 -613
rect 2589 -647 2623 -613
rect 2657 -647 2691 -613
rect 2725 -647 2759 -613
rect 2793 -647 2827 -613
rect 2861 -647 2895 -613
rect 2929 -647 2963 -613
rect 2997 -647 3031 -613
rect 3065 -647 3099 -613
rect 3133 -647 3167 -613
rect 3201 -647 3235 -613
rect 3269 -647 3303 -613
rect 3337 -647 3371 -613
rect 3405 -647 3439 -613
rect 3473 -647 3507 -613
rect 3541 -647 3575 -613
rect 3609 -647 3643 -613
rect 3677 -647 3711 -613
rect 3745 -647 3779 -613
rect 3813 -647 3847 -613
rect 3881 -647 3915 -613
rect 3949 -647 3983 -613
rect 4017 -647 4051 -613
rect 4085 -647 4119 -613
rect 4153 -647 4187 -613
rect 4221 -647 4255 -613
rect 4289 -647 4323 -613
rect 4357 -647 4391 -613
rect 4425 -647 4459 -613
rect 4493 -647 4527 -613
rect 4561 -647 4595 -613
rect 4629 -647 4663 -613
rect 4697 -647 4731 -613
rect 4765 -647 4799 -613
rect 4833 -647 4867 -613
rect 4901 -647 4935 -613
rect 4969 -647 5003 -613
rect 5037 -647 5071 -613
rect 5105 -647 5139 -613
rect 5173 -647 5207 -613
rect 5241 -647 5275 -613
rect 5309 -647 5343 -613
rect 5377 -647 5411 -613
rect 5445 -647 5479 -613
rect 5513 -647 5547 -613
rect 5581 -647 5615 -613
rect 5649 -647 5683 -613
rect 5717 -647 5751 -613
rect 5785 -647 5819 -613
rect 5853 -647 5887 -613
rect 5921 -647 5955 -613
rect 5989 -647 6023 -613
rect 6057 -647 6091 -613
rect 6125 -647 6159 -613
rect 6193 -647 6227 -613
rect 6261 -647 6295 -613
rect 6329 -647 6363 -613
rect 6397 -647 6431 -613
rect 6465 -647 6499 -613
rect 6533 -647 6567 -613
rect 6601 -647 6635 -613
rect 6669 -647 6757 -613
<< metal1 >>
rect -520 4930 -160 5260
rect -520 4870 6300 4930
rect -140 4670 -80 4870
rect 440 4670 500 4870
rect 1020 4670 1080 4870
rect 1600 4670 1660 4870
rect 2180 4670 2240 4870
rect 2760 4670 2820 4870
rect 3340 4670 3400 4870
rect 3920 4670 3980 4870
rect 4500 4670 4560 4870
rect 5080 4670 5140 4870
rect 5660 4670 5720 4870
rect 6240 4670 6300 4870
rect -520 4430 -80 4670
rect 60 4610 500 4670
rect 640 4610 1080 4670
rect 1220 4610 1660 4670
rect 1800 4610 1940 4670
rect 2010 4610 2240 4670
rect 2380 4610 2820 4670
rect 2960 4610 3400 4670
rect 3540 4610 3980 4670
rect 4120 4610 4560 4670
rect 4700 4610 5140 4670
rect 5280 4610 5720 4670
rect 1790 4576 2140 4580
rect 1790 4524 1814 4576
rect 1866 4524 1939 4576
rect 1991 4524 2064 4576
rect 2116 4524 2140 4576
rect 40 4486 390 4490
rect 40 4434 64 4486
rect 116 4434 189 4486
rect 241 4434 314 4486
rect 366 4434 390 4486
rect 40 4430 390 4434
rect 630 4486 980 4490
rect 630 4434 654 4486
rect 706 4434 779 4486
rect 831 4434 904 4486
rect 956 4434 980 4486
rect 630 4430 980 4434
rect 1210 4486 1560 4490
rect 1210 4434 1234 4486
rect 1286 4434 1359 4486
rect 1411 4434 1484 4486
rect 1536 4434 1560 4486
rect 1210 4430 1560 4434
rect 1790 4430 2140 4524
rect 2370 4576 2720 4580
rect 2370 4524 2394 4576
rect 2446 4524 2519 4576
rect 2571 4524 2644 4576
rect 2696 4524 2720 4576
rect 2370 4430 2720 4524
rect 4110 4576 4460 4580
rect 4110 4524 4134 4576
rect 4186 4524 4259 4576
rect 4311 4524 4384 4576
rect 4436 4524 4460 4576
rect 2950 4486 3300 4490
rect 2950 4434 2974 4486
rect 3026 4434 3099 4486
rect 3151 4434 3224 4486
rect 3276 4434 3300 4486
rect 2950 4430 3300 4434
rect 3530 4486 3880 4490
rect 3530 4434 3554 4486
rect 3606 4434 3679 4486
rect 3731 4434 3804 4486
rect 3856 4434 3880 4486
rect 3530 4430 3880 4434
rect 4110 4430 4460 4524
rect 4690 4576 5040 4580
rect 4690 4524 4714 4576
rect 4766 4524 4839 4576
rect 4891 4524 4964 4576
rect 5016 4524 5040 4576
rect 4690 4430 5040 4524
rect 5260 4576 5610 4580
rect 5260 4524 5284 4576
rect 5336 4524 5409 4576
rect 5461 4524 5534 4576
rect 5586 4524 5610 4576
rect 5260 4430 5610 4524
rect 5860 4430 6300 4670
rect -140 2430 -80 4430
rect -520 2060 -80 2430
rect 70 2426 360 2430
rect 70 2374 94 2426
rect 146 2374 189 2426
rect 241 2374 284 2426
rect 336 2374 360 2426
rect 70 2370 360 2374
rect 440 2340 500 4140
rect 650 2426 940 2430
rect 650 2374 674 2426
rect 726 2374 769 2426
rect 821 2374 864 2426
rect 916 2374 940 2426
rect 650 2370 940 2374
rect 1020 2340 1080 4140
rect 1230 2426 1520 2430
rect 1230 2374 1254 2426
rect 1306 2374 1349 2426
rect 1401 2374 1444 2426
rect 1496 2374 1520 2426
rect 1230 2370 1520 2374
rect 1600 2340 1660 4140
rect 2180 2430 2240 4140
rect 2760 2430 2820 4140
rect 1810 2426 2100 2430
rect 1810 2374 1834 2426
rect 1886 2374 1929 2426
rect 1981 2374 2024 2426
rect 2076 2374 2100 2426
rect 1810 2370 2100 2374
rect 2180 2370 2330 2430
rect 2390 2426 2680 2430
rect 2390 2374 2414 2426
rect 2466 2374 2509 2426
rect 2561 2374 2604 2426
rect 2656 2374 2680 2426
rect 2390 2370 2680 2374
rect 2760 2370 2910 2430
rect 2970 2426 3260 2430
rect 2970 2374 2994 2426
rect 3046 2374 3089 2426
rect 3141 2374 3184 2426
rect 3236 2374 3260 2426
rect 2970 2370 3260 2374
rect 390 2326 550 2340
rect 390 2274 404 2326
rect 456 2274 484 2326
rect 536 2274 550 2326
rect 390 2260 550 2274
rect 970 2326 1130 2340
rect 970 2274 984 2326
rect 1036 2274 1064 2326
rect 1116 2274 1130 2326
rect 970 2260 1130 2274
rect 1550 2326 1710 2340
rect 1550 2274 1564 2326
rect 1616 2274 1644 2326
rect 1696 2274 1710 2326
rect 1550 2260 1710 2274
rect 2080 2326 2240 2340
rect 2080 2274 2094 2326
rect 2146 2274 2174 2326
rect 2226 2274 2240 2326
rect 2080 2260 2240 2274
rect 390 2216 550 2230
rect 390 2164 404 2216
rect 456 2164 484 2216
rect 536 2164 550 2216
rect 390 2150 550 2164
rect 970 2216 1130 2230
rect 970 2164 984 2216
rect 1036 2164 1064 2216
rect 1116 2164 1130 2216
rect 970 2150 1130 2164
rect 1550 2216 1710 2230
rect 1550 2164 1564 2216
rect 1616 2164 1644 2216
rect 1696 2164 1710 2216
rect 1550 2150 1710 2164
rect -140 60 -80 2060
rect -520 -180 -80 60
rect -140 -380 -80 -180
rect -520 -384 -80 -380
rect -520 -436 -486 -384
rect -434 -436 -386 -384
rect -334 -436 -286 -384
rect -234 -436 -80 -384
rect -520 -440 -80 -436
rect -50 2060 360 2120
rect -50 -470 10 2060
rect 440 350 500 2150
rect 530 2060 940 2120
rect 70 56 360 60
rect 70 4 94 56
rect 146 4 189 56
rect 241 4 284 56
rect 336 4 360 56
rect 70 0 360 4
rect 60 -180 500 -120
rect 440 -380 500 -180
rect 60 -384 500 -380
rect 60 -436 94 -384
rect 146 -436 194 -384
rect 246 -436 294 -384
rect 346 -436 500 -384
rect 60 -440 500 -436
rect 530 -470 590 2060
rect 1020 350 1080 2150
rect 1110 2060 1520 2120
rect 650 56 940 60
rect 650 4 674 56
rect 726 4 769 56
rect 821 4 864 56
rect 916 4 940 56
rect 650 0 940 4
rect 640 -180 1080 -120
rect 1020 -380 1080 -180
rect 640 -384 1080 -380
rect 640 -436 674 -384
rect 726 -436 774 -384
rect 826 -436 874 -384
rect 926 -436 1080 -384
rect 640 -440 1080 -436
rect 1110 -470 1170 2060
rect 1600 350 1660 2150
rect 1690 2060 2100 2120
rect 1230 56 1520 60
rect 1230 4 1254 56
rect 1306 4 1349 56
rect 1401 4 1444 56
rect 1496 4 1520 56
rect 1230 0 1520 4
rect 1690 -30 1750 2060
rect 2180 350 2240 2260
rect 2270 2230 2330 2370
rect 2660 2326 2820 2340
rect 2660 2274 2674 2326
rect 2726 2274 2754 2326
rect 2806 2274 2820 2326
rect 2660 2260 2820 2274
rect 2270 2216 2430 2230
rect 2270 2164 2284 2216
rect 2336 2164 2364 2216
rect 2416 2164 2430 2216
rect 2270 2150 2430 2164
rect 2270 2060 2680 2120
rect 1810 56 2100 60
rect 1810 4 1834 56
rect 1886 4 1929 56
rect 1981 4 2024 56
rect 2076 4 2100 56
rect 1810 0 2100 4
rect 2270 -30 2330 2060
rect 2760 350 2820 2260
rect 2850 2230 2910 2370
rect 3340 2340 3400 4140
rect 3550 2426 3840 2430
rect 3550 2374 3574 2426
rect 3626 2374 3669 2426
rect 3721 2374 3764 2426
rect 3816 2374 3840 2426
rect 3550 2370 3840 2374
rect 3920 2340 3980 4140
rect 4500 2430 4560 4140
rect 5080 2430 5140 4140
rect 5660 2430 5720 4140
rect 6240 2430 6300 4430
rect 4130 2426 4420 2430
rect 4130 2374 4154 2426
rect 4206 2374 4249 2426
rect 4301 2374 4344 2426
rect 4396 2374 4420 2426
rect 4130 2370 4420 2374
rect 4500 2370 4650 2430
rect 4710 2426 5000 2430
rect 4710 2374 4734 2426
rect 4786 2374 4829 2426
rect 4881 2374 4924 2426
rect 4976 2374 5000 2426
rect 4710 2370 5000 2374
rect 5080 2370 5230 2430
rect 5290 2426 5580 2430
rect 5290 2374 5314 2426
rect 5366 2374 5409 2426
rect 5461 2374 5504 2426
rect 5556 2374 5580 2426
rect 5290 2370 5580 2374
rect 5660 2370 5810 2430
rect 5860 2370 6300 2430
rect 3290 2326 3450 2340
rect 3290 2274 3304 2326
rect 3356 2274 3384 2326
rect 3436 2274 3450 2326
rect 3290 2260 3450 2274
rect 3870 2326 4030 2340
rect 3870 2274 3884 2326
rect 3936 2274 3964 2326
rect 4016 2274 4030 2326
rect 3870 2260 4030 2274
rect 4400 2326 4560 2340
rect 4400 2274 4414 2326
rect 4466 2274 4494 2326
rect 4546 2274 4560 2326
rect 4400 2260 4560 2274
rect 2850 2216 3010 2230
rect 2850 2164 2864 2216
rect 2916 2164 2944 2216
rect 2996 2164 3010 2216
rect 2850 2150 3010 2164
rect 3290 2216 3450 2230
rect 3290 2164 3304 2216
rect 3356 2164 3384 2216
rect 3436 2164 3450 2216
rect 3290 2150 3450 2164
rect 3870 2216 4030 2230
rect 3870 2164 3884 2216
rect 3936 2164 3964 2216
rect 4016 2164 4030 2216
rect 3870 2150 4030 2164
rect 2850 2060 3260 2120
rect 2390 56 2680 60
rect 2390 4 2414 56
rect 2466 4 2509 56
rect 2561 4 2604 56
rect 2656 4 2680 56
rect 2390 0 2680 4
rect 1640 -34 1800 -30
rect 1640 -86 1654 -34
rect 1706 -86 1734 -34
rect 1786 -86 1800 -34
rect 1640 -90 1800 -86
rect 2220 -34 2380 -30
rect 2220 -86 2234 -34
rect 2286 -86 2314 -34
rect 2366 -86 2380 -34
rect 2220 -90 2380 -86
rect 1220 -180 1660 -120
rect 1800 -180 2240 -120
rect 2380 -180 2820 -120
rect 1600 -380 1660 -180
rect 2180 -380 2240 -180
rect 2760 -380 2820 -180
rect 1220 -384 1660 -380
rect 1220 -436 1254 -384
rect 1306 -436 1354 -384
rect 1406 -436 1454 -384
rect 1506 -436 1660 -384
rect 1220 -440 1660 -436
rect 1800 -384 2240 -380
rect 1800 -436 1834 -384
rect 1886 -436 1934 -384
rect 1986 -436 2034 -384
rect 2086 -436 2240 -384
rect 1800 -440 2240 -436
rect 2380 -384 2820 -380
rect 2380 -436 2414 -384
rect 2466 -436 2514 -384
rect 2566 -436 2614 -384
rect 2666 -436 2820 -384
rect 2380 -440 2820 -436
rect 2850 -470 2910 2060
rect 3340 350 3400 2150
rect 3430 2060 3840 2120
rect 2970 56 3260 60
rect 2970 4 2994 56
rect 3046 4 3089 56
rect 3141 4 3184 56
rect 3236 4 3260 56
rect 2970 0 3260 4
rect 2960 -180 3400 -120
rect 3340 -380 3400 -180
rect 2960 -384 3400 -380
rect 2960 -436 2994 -384
rect 3046 -436 3094 -384
rect 3146 -436 3194 -384
rect 3246 -436 3400 -384
rect 2960 -440 3400 -436
rect 3430 -470 3490 2060
rect 3920 350 3980 2150
rect 4010 2060 4420 2120
rect 3550 56 3840 60
rect 3550 4 3574 56
rect 3626 4 3669 56
rect 3721 4 3764 56
rect 3816 4 3840 56
rect 3550 0 3840 4
rect 4010 -30 4070 2060
rect 4500 350 4560 2260
rect 4590 2230 4650 2370
rect 4980 2326 5140 2340
rect 4980 2274 4994 2326
rect 5046 2274 5074 2326
rect 5126 2274 5140 2326
rect 4980 2260 5140 2274
rect 4590 2216 4750 2230
rect 4590 2164 4604 2216
rect 4656 2164 4684 2216
rect 4736 2164 4750 2216
rect 4590 2150 4750 2164
rect 4590 2060 5000 2120
rect 4130 56 4420 60
rect 4130 4 4154 56
rect 4206 4 4249 56
rect 4301 4 4344 56
rect 4396 4 4420 56
rect 4130 0 4420 4
rect 4590 -30 4650 2060
rect 5080 350 5140 2260
rect 5170 2230 5230 2370
rect 5560 2326 5720 2340
rect 5560 2274 5574 2326
rect 5626 2274 5654 2326
rect 5706 2274 5720 2326
rect 5560 2260 5720 2274
rect 5170 2216 5330 2230
rect 5170 2164 5184 2216
rect 5236 2164 5264 2216
rect 5316 2164 5330 2216
rect 5170 2150 5330 2164
rect 5170 2060 5580 2120
rect 4710 56 5000 60
rect 4710 4 4734 56
rect 4786 4 4829 56
rect 4881 4 4924 56
rect 4976 4 5000 56
rect 4710 0 5000 4
rect 5170 -30 5230 2060
rect 5660 350 5720 2260
rect 5750 2230 5810 2370
rect 5750 2216 5910 2230
rect 5750 2164 5764 2216
rect 5816 2164 5844 2216
rect 5896 2164 5910 2216
rect 5750 2150 5910 2164
rect 5950 2120 6300 2370
rect 5860 2060 6300 2120
rect 6240 60 6300 2060
rect 5290 56 5580 60
rect 5290 4 5314 56
rect 5366 4 5409 56
rect 5461 4 5504 56
rect 5556 4 5580 56
rect 5290 0 5580 4
rect 3960 -34 4120 -30
rect 3960 -86 3974 -34
rect 4026 -86 4054 -34
rect 4106 -86 4120 -34
rect 3960 -90 4120 -86
rect 4540 -34 4700 -30
rect 4540 -86 4554 -34
rect 4606 -86 4634 -34
rect 4686 -86 4700 -34
rect 4540 -90 4700 -86
rect 5120 -34 5280 -30
rect 5120 -86 5134 -34
rect 5186 -86 5214 -34
rect 5266 -86 5280 -34
rect 5120 -90 5280 -86
rect 3540 -180 3980 -120
rect 4120 -180 4560 -120
rect 4700 -180 5140 -120
rect 5280 -180 5720 -120
rect 5860 -180 6300 60
rect 3920 -380 3980 -180
rect 4500 -380 4560 -180
rect 5080 -380 5140 -180
rect 5660 -380 5720 -180
rect 6240 -380 6300 -180
rect 3540 -384 3980 -380
rect 3540 -436 3574 -384
rect 3626 -436 3674 -384
rect 3726 -436 3774 -384
rect 3826 -436 3980 -384
rect 3540 -440 3980 -436
rect 4120 -384 4560 -380
rect 4120 -436 4154 -384
rect 4206 -436 4254 -384
rect 4306 -436 4354 -384
rect 4406 -436 4560 -384
rect 4120 -440 4560 -436
rect 4700 -384 5140 -380
rect 4700 -436 4734 -384
rect 4786 -436 4834 -384
rect 4886 -436 4934 -384
rect 4986 -436 5140 -384
rect 4700 -440 5140 -436
rect 5280 -384 5720 -380
rect 5280 -436 5304 -384
rect 5356 -436 5404 -384
rect 5456 -436 5504 -384
rect 5556 -436 5720 -384
rect 5280 -440 5720 -436
rect 5860 -384 6300 -380
rect 5860 -436 5884 -384
rect 5936 -436 5984 -384
rect 6036 -436 6084 -384
rect 6136 -436 6300 -384
rect 5860 -440 6300 -436
rect -100 -474 60 -470
rect -100 -526 -86 -474
rect -34 -526 -6 -474
rect 46 -526 60 -474
rect -100 -530 60 -526
rect 480 -474 640 -470
rect 480 -526 494 -474
rect 546 -526 574 -474
rect 626 -526 640 -474
rect 480 -530 640 -526
rect 1060 -474 1220 -470
rect 1060 -526 1074 -474
rect 1126 -526 1154 -474
rect 1206 -526 1220 -474
rect 1060 -530 1220 -526
rect 2800 -474 2960 -470
rect 2800 -526 2814 -474
rect 2866 -526 2894 -474
rect 2946 -526 2960 -474
rect 2800 -530 2960 -526
rect 3380 -474 3540 -470
rect 3380 -526 3394 -474
rect 3446 -526 3474 -474
rect 3526 -526 3540 -474
rect 3380 -530 3540 -526
<< via1 >>
rect 1814 4524 1866 4576
rect 1939 4524 1991 4576
rect 2064 4524 2116 4576
rect 64 4434 116 4486
rect 189 4434 241 4486
rect 314 4434 366 4486
rect 654 4434 706 4486
rect 779 4434 831 4486
rect 904 4434 956 4486
rect 1234 4434 1286 4486
rect 1359 4434 1411 4486
rect 1484 4434 1536 4486
rect 2394 4524 2446 4576
rect 2519 4524 2571 4576
rect 2644 4524 2696 4576
rect 4134 4524 4186 4576
rect 4259 4524 4311 4576
rect 4384 4524 4436 4576
rect 2974 4434 3026 4486
rect 3099 4434 3151 4486
rect 3224 4434 3276 4486
rect 3554 4434 3606 4486
rect 3679 4434 3731 4486
rect 3804 4434 3856 4486
rect 4714 4524 4766 4576
rect 4839 4524 4891 4576
rect 4964 4524 5016 4576
rect 5284 4524 5336 4576
rect 5409 4524 5461 4576
rect 5534 4524 5586 4576
rect 94 2374 146 2426
rect 189 2374 241 2426
rect 284 2374 336 2426
rect 674 2374 726 2426
rect 769 2374 821 2426
rect 864 2374 916 2426
rect 1254 2374 1306 2426
rect 1349 2374 1401 2426
rect 1444 2374 1496 2426
rect 1834 2374 1886 2426
rect 1929 2374 1981 2426
rect 2024 2374 2076 2426
rect 2414 2374 2466 2426
rect 2509 2374 2561 2426
rect 2604 2374 2656 2426
rect 2994 2374 3046 2426
rect 3089 2374 3141 2426
rect 3184 2374 3236 2426
rect 404 2274 456 2326
rect 484 2274 536 2326
rect 984 2274 1036 2326
rect 1064 2274 1116 2326
rect 1564 2274 1616 2326
rect 1644 2274 1696 2326
rect 2094 2274 2146 2326
rect 2174 2274 2226 2326
rect 404 2164 456 2216
rect 484 2164 536 2216
rect 984 2164 1036 2216
rect 1064 2164 1116 2216
rect 1564 2164 1616 2216
rect 1644 2164 1696 2216
rect -486 -436 -434 -384
rect -386 -436 -334 -384
rect -286 -436 -234 -384
rect 94 4 146 56
rect 189 4 241 56
rect 284 4 336 56
rect 94 -436 146 -384
rect 194 -436 246 -384
rect 294 -436 346 -384
rect 674 4 726 56
rect 769 4 821 56
rect 864 4 916 56
rect 674 -436 726 -384
rect 774 -436 826 -384
rect 874 -436 926 -384
rect 1254 4 1306 56
rect 1349 4 1401 56
rect 1444 4 1496 56
rect 2674 2274 2726 2326
rect 2754 2274 2806 2326
rect 2284 2164 2336 2216
rect 2364 2164 2416 2216
rect 1834 4 1886 56
rect 1929 4 1981 56
rect 2024 4 2076 56
rect 3574 2374 3626 2426
rect 3669 2374 3721 2426
rect 3764 2374 3816 2426
rect 4154 2374 4206 2426
rect 4249 2374 4301 2426
rect 4344 2374 4396 2426
rect 4734 2374 4786 2426
rect 4829 2374 4881 2426
rect 4924 2374 4976 2426
rect 5314 2374 5366 2426
rect 5409 2374 5461 2426
rect 5504 2374 5556 2426
rect 3304 2274 3356 2326
rect 3384 2274 3436 2326
rect 3884 2274 3936 2326
rect 3964 2274 4016 2326
rect 4414 2274 4466 2326
rect 4494 2274 4546 2326
rect 2864 2164 2916 2216
rect 2944 2164 2996 2216
rect 3304 2164 3356 2216
rect 3384 2164 3436 2216
rect 3884 2164 3936 2216
rect 3964 2164 4016 2216
rect 2414 4 2466 56
rect 2509 4 2561 56
rect 2604 4 2656 56
rect 1654 -86 1706 -34
rect 1734 -86 1786 -34
rect 2234 -86 2286 -34
rect 2314 -86 2366 -34
rect 1254 -436 1306 -384
rect 1354 -436 1406 -384
rect 1454 -436 1506 -384
rect 1834 -436 1886 -384
rect 1934 -436 1986 -384
rect 2034 -436 2086 -384
rect 2414 -436 2466 -384
rect 2514 -436 2566 -384
rect 2614 -436 2666 -384
rect 2994 4 3046 56
rect 3089 4 3141 56
rect 3184 4 3236 56
rect 2994 -436 3046 -384
rect 3094 -436 3146 -384
rect 3194 -436 3246 -384
rect 3574 4 3626 56
rect 3669 4 3721 56
rect 3764 4 3816 56
rect 4994 2274 5046 2326
rect 5074 2274 5126 2326
rect 4604 2164 4656 2216
rect 4684 2164 4736 2216
rect 4154 4 4206 56
rect 4249 4 4301 56
rect 4344 4 4396 56
rect 5574 2274 5626 2326
rect 5654 2274 5706 2326
rect 5184 2164 5236 2216
rect 5264 2164 5316 2216
rect 4734 4 4786 56
rect 4829 4 4881 56
rect 4924 4 4976 56
rect 5764 2164 5816 2216
rect 5844 2164 5896 2216
rect 5314 4 5366 56
rect 5409 4 5461 56
rect 5504 4 5556 56
rect 3974 -86 4026 -34
rect 4054 -86 4106 -34
rect 4554 -86 4606 -34
rect 4634 -86 4686 -34
rect 5134 -86 5186 -34
rect 5214 -86 5266 -34
rect 3574 -436 3626 -384
rect 3674 -436 3726 -384
rect 3774 -436 3826 -384
rect 4154 -436 4206 -384
rect 4254 -436 4306 -384
rect 4354 -436 4406 -384
rect 4734 -436 4786 -384
rect 4834 -436 4886 -384
rect 4934 -436 4986 -384
rect 5304 -436 5356 -384
rect 5404 -436 5456 -384
rect 5504 -436 5556 -384
rect 5884 -436 5936 -384
rect 5984 -436 6036 -384
rect 6084 -436 6136 -384
rect -86 -526 -34 -474
rect -6 -526 46 -474
rect 494 -526 546 -474
rect 574 -526 626 -474
rect 1074 -526 1126 -474
rect 1154 -526 1206 -474
rect 2814 -526 2866 -474
rect 2894 -526 2946 -474
rect 3394 -526 3446 -474
rect 3474 -526 3526 -474
<< metal2 >>
rect 1800 4763 1940 4800
rect 1800 4707 1842 4763
rect 1898 4707 1940 4763
rect 10 4548 150 4590
rect 1800 4580 1940 4707
rect 10 4492 52 4548
rect 108 4492 150 4548
rect 1790 4576 6680 4580
rect 1790 4524 1814 4576
rect 1866 4524 1939 4576
rect 1991 4524 2064 4576
rect 2116 4524 2394 4576
rect 2446 4524 2519 4576
rect 2571 4524 2644 4576
rect 2696 4524 4134 4576
rect 4186 4524 4259 4576
rect 4311 4524 4384 4576
rect 4436 4524 4714 4576
rect 4766 4524 4839 4576
rect 4891 4524 4964 4576
rect 5016 4524 5284 4576
rect 5336 4524 5409 4576
rect 5461 4524 5534 4576
rect 5586 4568 6680 4576
rect 5586 4524 6612 4568
rect 1790 4520 6612 4524
rect 10 4490 150 4492
rect 6600 4512 6612 4520
rect 6668 4512 6680 4568
rect 10 4486 6540 4490
rect 10 4434 64 4486
rect 116 4434 189 4486
rect 241 4434 314 4486
rect 366 4434 654 4486
rect 706 4434 779 4486
rect 831 4434 904 4486
rect 956 4434 1234 4486
rect 1286 4434 1359 4486
rect 1411 4434 1484 4486
rect 1536 4434 2974 4486
rect 3026 4434 3099 4486
rect 3151 4434 3224 4486
rect 3276 4434 3554 4486
rect 3606 4434 3679 4486
rect 3731 4434 3804 4486
rect 3856 4478 6540 4486
rect 3856 4434 6472 4478
rect 10 4430 6472 4434
rect 6460 4422 6472 4430
rect 6528 4422 6540 4478
rect 6460 4388 6540 4422
rect 6600 4478 6680 4512
rect 6600 4422 6612 4478
rect 6668 4422 6680 4478
rect 6600 4410 6680 4422
rect 6460 4332 6472 4388
rect 6528 4332 6540 4388
rect 6460 4320 6540 4332
rect -1010 2418 -910 2440
rect -1010 2362 -988 2418
rect -932 2362 -910 2418
rect 30 2426 6400 2430
rect 30 2374 94 2426
rect 146 2374 189 2426
rect 241 2374 284 2426
rect 336 2374 674 2426
rect 726 2374 769 2426
rect 821 2374 864 2426
rect 916 2374 1254 2426
rect 1306 2374 1349 2426
rect 1401 2374 1444 2426
rect 1496 2374 1834 2426
rect 1886 2374 1929 2426
rect 1981 2374 2024 2426
rect 2076 2374 2414 2426
rect 2466 2374 2509 2426
rect 2561 2374 2604 2426
rect 2656 2374 2994 2426
rect 3046 2374 3089 2426
rect 3141 2374 3184 2426
rect 3236 2374 3574 2426
rect 3626 2374 3669 2426
rect 3721 2374 3764 2426
rect 3816 2374 4154 2426
rect 4206 2374 4249 2426
rect 4301 2374 4344 2426
rect 4396 2374 4734 2426
rect 4786 2374 4829 2426
rect 4881 2374 4924 2426
rect 4976 2374 5314 2426
rect 5366 2374 5409 2426
rect 5461 2374 5504 2426
rect 5556 2418 6400 2426
rect 5556 2374 6332 2418
rect 30 2370 6332 2374
rect -1010 2340 -910 2362
rect 6320 2362 6332 2370
rect 6388 2362 6400 2418
rect -1000 2326 5720 2340
rect -1000 2274 404 2326
rect 456 2274 484 2326
rect 536 2274 984 2326
rect 1036 2274 1064 2326
rect 1116 2274 1564 2326
rect 1616 2274 1644 2326
rect 1696 2274 2094 2326
rect 2146 2274 2174 2326
rect 2226 2274 2674 2326
rect 2726 2274 2754 2326
rect 2806 2274 3304 2326
rect 3356 2274 3384 2326
rect 3436 2274 3884 2326
rect 3936 2274 3964 2326
rect 4016 2274 4414 2326
rect 4466 2274 4494 2326
rect 4546 2274 4994 2326
rect 5046 2274 5074 2326
rect 5126 2274 5574 2326
rect 5626 2274 5654 2326
rect 5706 2274 5720 2326
rect -1000 2260 5720 2274
rect 6320 2328 6400 2362
rect 6320 2272 6332 2328
rect 6388 2272 6400 2328
rect 6320 2260 6400 2272
rect -1000 2216 5910 2230
rect -1000 2164 404 2216
rect 456 2164 484 2216
rect 536 2164 984 2216
rect 1036 2164 1064 2216
rect 1116 2164 1564 2216
rect 1616 2164 1644 2216
rect 1696 2164 2284 2216
rect 2336 2164 2364 2216
rect 2416 2164 2864 2216
rect 2916 2164 2944 2216
rect 2996 2164 3304 2216
rect 3356 2164 3384 2216
rect 3436 2164 3884 2216
rect 3936 2164 3964 2216
rect 4016 2164 4604 2216
rect 4656 2164 4684 2216
rect 4736 2164 5184 2216
rect 5236 2164 5264 2216
rect 5316 2164 5764 2216
rect 5816 2164 5844 2216
rect 5896 2164 5910 2216
rect -1000 2150 5910 2164
rect -1010 2128 -910 2150
rect -1010 2072 -988 2128
rect -932 2072 -910 2128
rect -1010 2050 -910 2072
rect 6320 158 6400 170
rect 6320 102 6332 158
rect 6388 102 6400 158
rect 6320 70 6400 102
rect 6810 70 6910 90
rect 6320 68 6910 70
rect 6320 60 6332 68
rect 50 56 6332 60
rect 50 4 94 56
rect 146 4 189 56
rect 241 4 284 56
rect 336 4 674 56
rect 726 4 769 56
rect 821 4 864 56
rect 916 4 1254 56
rect 1306 4 1349 56
rect 1401 4 1444 56
rect 1496 4 1834 56
rect 1886 4 1929 56
rect 1981 4 2024 56
rect 2076 4 2414 56
rect 2466 4 2509 56
rect 2561 4 2604 56
rect 2656 4 2994 56
rect 3046 4 3089 56
rect 3141 4 3184 56
rect 3236 4 3574 56
rect 3626 4 3669 56
rect 3721 4 3764 56
rect 3816 4 4154 56
rect 4206 4 4249 56
rect 4301 4 4344 56
rect 4396 4 4734 56
rect 4786 4 4829 56
rect 4881 4 4924 56
rect 4976 4 5314 56
rect 5366 4 5409 56
rect 5461 4 5504 56
rect 5556 12 6332 56
rect 6388 63 6910 68
rect 6388 12 6832 63
rect 5556 7 6832 12
rect 6888 7 6910 63
rect 5556 4 6910 7
rect 50 0 6910 4
rect 6810 -20 6910 0
rect 1640 -34 6540 -30
rect 1640 -86 1654 -34
rect 1706 -86 1734 -34
rect 1786 -86 2234 -34
rect 2286 -86 2314 -34
rect 2366 -86 3974 -34
rect 4026 -86 4054 -34
rect 4106 -86 4554 -34
rect 4606 -86 4634 -34
rect 4686 -86 5134 -34
rect 5186 -86 5214 -34
rect 5266 -42 6540 -34
rect 5266 -86 6472 -42
rect 1640 -90 6472 -86
rect 6460 -98 6472 -90
rect 6528 -98 6540 -42
rect 6460 -132 6540 -98
rect 6460 -188 6472 -132
rect 6528 -188 6540 -132
rect 6460 -200 6540 -188
rect 6600 -372 6680 -360
rect -520 -384 6170 -380
rect -520 -436 -486 -384
rect -434 -436 -386 -384
rect -334 -436 -286 -384
rect -234 -436 94 -384
rect 146 -436 194 -384
rect 246 -436 294 -384
rect 346 -436 674 -384
rect 726 -436 774 -384
rect 826 -436 874 -384
rect 926 -436 1254 -384
rect 1306 -436 1354 -384
rect 1406 -436 1454 -384
rect 1506 -436 1834 -384
rect 1886 -436 1934 -384
rect 1986 -436 2034 -384
rect 2086 -436 2414 -384
rect 2466 -436 2514 -384
rect 2566 -436 2614 -384
rect 2666 -436 2994 -384
rect 3046 -436 3094 -384
rect 3146 -436 3194 -384
rect 3246 -436 3574 -384
rect 3626 -436 3674 -384
rect 3726 -436 3774 -384
rect 3826 -436 4154 -384
rect 4206 -436 4254 -384
rect 4306 -436 4354 -384
rect 4406 -436 4734 -384
rect 4786 -436 4834 -384
rect 4886 -436 4934 -384
rect 4986 -436 5304 -384
rect 5356 -436 5404 -384
rect 5456 -436 5504 -384
rect 5556 -436 5884 -384
rect 5936 -436 5984 -384
rect 6036 -436 6084 -384
rect 6136 -436 6170 -384
rect -520 -440 6170 -436
rect 6600 -428 6612 -372
rect 6668 -428 6680 -372
rect 6600 -462 6680 -428
rect 6600 -470 6612 -462
rect -100 -474 6612 -470
rect -100 -526 -86 -474
rect -34 -526 -6 -474
rect 46 -526 494 -474
rect 546 -526 574 -474
rect 626 -526 1074 -474
rect 1126 -526 1154 -474
rect 1206 -526 2814 -474
rect 2866 -526 2894 -474
rect 2946 -526 3394 -474
rect 3446 -526 3474 -474
rect 3526 -518 6612 -474
rect 6668 -518 6680 -462
rect 3526 -526 6680 -518
rect -100 -530 6680 -526
<< via2 >>
rect 1842 4707 1898 4763
rect 52 4492 108 4548
rect 6612 4512 6668 4568
rect 6472 4422 6528 4478
rect 6612 4422 6668 4478
rect 6472 4332 6528 4388
rect -988 2362 -932 2418
rect 6332 2362 6388 2418
rect 6332 2272 6388 2328
rect -988 2072 -932 2128
rect 6332 102 6388 158
rect 6332 12 6388 68
rect 6832 7 6888 63
rect 6472 -98 6528 -42
rect 6472 -188 6528 -132
rect 6612 -428 6668 -372
rect 6612 -518 6668 -462
<< metal3 >>
rect 10 4548 150 5260
rect 1800 4763 1940 5260
rect 1800 4707 1842 4763
rect 1898 4707 1940 4763
rect 1800 4668 1940 4707
rect 10 4492 52 4548
rect 108 4492 150 4548
rect 10 4490 150 4492
rect 6600 4568 6680 4580
rect 6600 4512 6612 4568
rect 6668 4512 6680 4568
rect 10 4410 190 4490
rect 6460 4478 6540 4490
rect 6460 4422 6472 4478
rect 6528 4422 6540 4478
rect 6460 4388 6540 4422
rect 6460 4332 6472 4388
rect 6528 4332 6540 4388
rect -1010 2418 -910 2440
rect -1010 2362 -988 2418
rect -932 2362 -910 2418
rect -1010 2340 -910 2362
rect 6320 2418 6400 2430
rect 6320 2362 6332 2418
rect 6388 2362 6400 2418
rect 6320 2328 6400 2362
rect 6320 2272 6332 2328
rect 6388 2272 6400 2328
rect -1010 2128 -910 2150
rect -1010 2072 -988 2128
rect -932 2072 -910 2128
rect -1010 2050 -910 2072
rect 6320 158 6400 2272
rect 6320 102 6332 158
rect 6388 102 6400 158
rect 6320 68 6400 102
rect 6320 12 6332 68
rect 6388 12 6400 68
rect 6320 0 6400 12
rect 6460 -42 6540 4332
rect 6460 -98 6472 -42
rect 6528 -98 6540 -42
rect 6460 -132 6540 -98
rect 6460 -188 6472 -132
rect 6528 -188 6540 -132
rect 6460 -200 6540 -188
rect 6600 4478 6680 4512
rect 6600 4422 6612 4478
rect 6668 4422 6680 4478
rect 6600 -372 6680 4422
rect 6810 63 6910 90
rect 6810 7 6832 63
rect 6888 7 6910 63
rect 6810 -20 6910 7
rect 6600 -428 6612 -372
rect 6668 -428 6680 -372
rect 6600 -462 6680 -428
rect 6600 -518 6612 -462
rect 6668 -518 6680 -462
rect 6600 -530 6680 -518
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_0
timestamp 1757161594
transform 0 1 827 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_2
timestamp 1757161594
transform 0 1 1407 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_3
timestamp 1757161594
transform 0 1 1987 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_4
timestamp 1757161594
transform 0 1 2567 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_5
timestamp 1757161594
transform 0 1 3147 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_6
timestamp 1757161594
transform 0 1 3727 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_7
timestamp 1757161594
transform 0 1 4307 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_8
timestamp 1757161594
transform 0 1 4887 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_9
timestamp 1757161594
transform 0 1 5467 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_10
timestamp 1757161594
transform 0 1 6047 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_11
timestamp 1757161594
transform 0 1 -333 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_12
timestamp 1757161594
transform 0 1 -333 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_13
timestamp 1757161594
transform 0 1 827 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_14
timestamp 1757161594
transform 0 1 2567 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_15
timestamp 1757161594
transform 0 1 3147 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_16
timestamp 1757161594
transform 0 1 1407 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_17
timestamp 1757161594
transform 0 1 1987 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_18
timestamp 1757161594
transform 0 1 4887 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_19
timestamp 1757161594
transform 0 1 5467 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_20
timestamp 1757161594
transform 0 1 3727 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_21
timestamp 1757161594
transform 0 1 4307 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_22
timestamp 1757161594
transform 0 1 6047 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_24
timestamp 1757161594
transform 0 1 247 -1 0 -282
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_ND6TEZ  sky130_fd_pr__nfet_01v8_lvt_ND6TEZ_25
timestamp 1757161594
transform 0 1 247 -1 0 4768
box -184 -257 184 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_0
timestamp 1757161594
transform 0 1 5467 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_1
timestamp 1757161594
transform 0 1 3147 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_2
timestamp 1757161594
transform 0 1 3727 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_3
timestamp 1757161594
transform 0 1 4307 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_4
timestamp 1757161594
transform 0 1 4887 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_5
timestamp 1757161594
transform 0 1 2567 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_6
timestamp 1757161594
transform 0 1 1987 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_7
timestamp 1757161594
transform 0 1 1407 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_8
timestamp 1757161594
transform 0 1 827 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_9
timestamp 1757161594
transform 0 1 247 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_10
timestamp 1757161594
transform 0 1 6047 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_12
timestamp 1757161594
transform 0 1 5467 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_13
timestamp 1757161594
transform 0 1 4887 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_14
timestamp 1757161594
transform 0 1 4307 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_15
timestamp 1757161594
transform 0 1 3727 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_16
timestamp 1757161594
transform 0 1 3147 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_17
timestamp 1757161594
transform 0 1 2567 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_18
timestamp 1757161594
transform 0 1 1987 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_19
timestamp 1757161594
transform 0 1 1407 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_20
timestamp 1757161594
transform 0 1 827 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_21
timestamp 1757161594
transform 0 1 -333 -1 0 3428
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_22
timestamp 1757161594
transform 0 1 6047 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_24
timestamp 1757161594
transform 0 1 -333 -1 0 1058
box -1084 -257 1084 257
use sky130_fd_pr__nfet_01v8_lvt_VVFJJL  sky130_fd_pr__nfet_01v8_lvt_VVFJJL_25
timestamp 1757161594
transform 0 1 247 -1 0 3428
box -1084 -257 1084 257
<< labels >>
flabel metal2 s -1000 2340 -920 2420 0 FreeSans 1172 0 0 0 in-
port 1 nsew
flabel metal2 s -1000 2070 -920 2150 0 FreeSans 1172 0 0 0 in+
port 2 nsew
<< end >>
