magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -1196 -3076 2816 -2984
rect -1196 -5094 -1104 -3076
rect 2724 -5094 2816 -3076
rect -1196 -5226 2816 -5094
<< psubdiff >>
rect -1170 -3050 2790 -3010
rect -1170 -5120 -1130 -3050
rect 2750 -5120 2790 -3050
rect -1170 -5143 2790 -5120
rect -1170 -5177 -1111 -5143
rect -1077 -5177 -1043 -5143
rect -1009 -5177 -975 -5143
rect -941 -5177 -907 -5143
rect -873 -5177 -839 -5143
rect -805 -5177 -771 -5143
rect -737 -5177 -703 -5143
rect -669 -5177 -635 -5143
rect -601 -5177 -567 -5143
rect -533 -5177 -499 -5143
rect -465 -5177 -431 -5143
rect -397 -5177 -363 -5143
rect -329 -5177 -295 -5143
rect -261 -5177 -227 -5143
rect -193 -5177 -159 -5143
rect -125 -5177 -91 -5143
rect -57 -5177 -23 -5143
rect 11 -5177 45 -5143
rect 79 -5177 113 -5143
rect 147 -5177 181 -5143
rect 215 -5177 249 -5143
rect 283 -5177 317 -5143
rect 351 -5177 385 -5143
rect 419 -5177 453 -5143
rect 487 -5177 521 -5143
rect 555 -5177 589 -5143
rect 623 -5177 657 -5143
rect 691 -5177 725 -5143
rect 759 -5177 793 -5143
rect 827 -5177 861 -5143
rect 895 -5177 929 -5143
rect 963 -5177 997 -5143
rect 1031 -5177 1065 -5143
rect 1099 -5177 1133 -5143
rect 1167 -5177 1201 -5143
rect 1235 -5177 1269 -5143
rect 1303 -5177 1337 -5143
rect 1371 -5177 1405 -5143
rect 1439 -5177 1473 -5143
rect 1507 -5177 1541 -5143
rect 1575 -5177 1609 -5143
rect 1643 -5177 1677 -5143
rect 1711 -5177 1745 -5143
rect 1779 -5177 1813 -5143
rect 1847 -5177 1881 -5143
rect 1915 -5177 1949 -5143
rect 1983 -5177 2017 -5143
rect 2051 -5177 2085 -5143
rect 2119 -5177 2153 -5143
rect 2187 -5177 2221 -5143
rect 2255 -5177 2289 -5143
rect 2323 -5177 2357 -5143
rect 2391 -5177 2425 -5143
rect 2459 -5177 2493 -5143
rect 2527 -5177 2561 -5143
rect 2595 -5177 2629 -5143
rect 2663 -5177 2697 -5143
rect 2731 -5177 2790 -5143
rect -1170 -5200 2790 -5177
<< psubdiffcont >>
rect -1111 -5177 -1077 -5143
rect -1043 -5177 -1009 -5143
rect -975 -5177 -941 -5143
rect -907 -5177 -873 -5143
rect -839 -5177 -805 -5143
rect -771 -5177 -737 -5143
rect -703 -5177 -669 -5143
rect -635 -5177 -601 -5143
rect -567 -5177 -533 -5143
rect -499 -5177 -465 -5143
rect -431 -5177 -397 -5143
rect -363 -5177 -329 -5143
rect -295 -5177 -261 -5143
rect -227 -5177 -193 -5143
rect -159 -5177 -125 -5143
rect -91 -5177 -57 -5143
rect -23 -5177 11 -5143
rect 45 -5177 79 -5143
rect 113 -5177 147 -5143
rect 181 -5177 215 -5143
rect 249 -5177 283 -5143
rect 317 -5177 351 -5143
rect 385 -5177 419 -5143
rect 453 -5177 487 -5143
rect 521 -5177 555 -5143
rect 589 -5177 623 -5143
rect 657 -5177 691 -5143
rect 725 -5177 759 -5143
rect 793 -5177 827 -5143
rect 861 -5177 895 -5143
rect 929 -5177 963 -5143
rect 997 -5177 1031 -5143
rect 1065 -5177 1099 -5143
rect 1133 -5177 1167 -5143
rect 1201 -5177 1235 -5143
rect 1269 -5177 1303 -5143
rect 1337 -5177 1371 -5143
rect 1405 -5177 1439 -5143
rect 1473 -5177 1507 -5143
rect 1541 -5177 1575 -5143
rect 1609 -5177 1643 -5143
rect 1677 -5177 1711 -5143
rect 1745 -5177 1779 -5143
rect 1813 -5177 1847 -5143
rect 1881 -5177 1915 -5143
rect 1949 -5177 1983 -5143
rect 2017 -5177 2051 -5143
rect 2085 -5177 2119 -5143
rect 2153 -5177 2187 -5143
rect 2221 -5177 2255 -5143
rect 2289 -5177 2323 -5143
rect 2357 -5177 2391 -5143
rect 2425 -5177 2459 -5143
rect 2493 -5177 2527 -5143
rect 2561 -5177 2595 -5143
rect 2629 -5177 2663 -5143
rect 2697 -5177 2731 -5143
<< locali >>
rect -1170 -3050 2790 -3010
rect -1170 -5120 -1130 -3050
rect 2750 -5120 2790 -3050
rect -1170 -5143 2790 -5120
rect -1170 -5177 -1115 -5143
rect -1077 -5177 -1043 -5143
rect -1009 -5177 -975 -5143
rect -937 -5177 -907 -5143
rect -865 -5177 -839 -5143
rect -793 -5177 -771 -5143
rect -721 -5177 -703 -5143
rect -649 -5177 -635 -5143
rect -577 -5177 -567 -5143
rect -505 -5177 -499 -5143
rect -433 -5177 -431 -5143
rect -397 -5177 -395 -5143
rect -329 -5177 -323 -5143
rect -261 -5177 -251 -5143
rect -193 -5177 -179 -5143
rect -125 -5177 -107 -5143
rect -57 -5177 -35 -5143
rect 11 -5177 37 -5143
rect 79 -5177 109 -5143
rect 147 -5177 181 -5143
rect 215 -5177 249 -5143
rect 287 -5177 317 -5143
rect 359 -5177 385 -5143
rect 431 -5177 453 -5143
rect 503 -5177 521 -5143
rect 575 -5177 589 -5143
rect 647 -5177 657 -5143
rect 719 -5177 725 -5143
rect 791 -5177 793 -5143
rect 827 -5177 829 -5143
rect 895 -5177 901 -5143
rect 963 -5177 973 -5143
rect 1031 -5177 1045 -5143
rect 1099 -5177 1117 -5143
rect 1167 -5177 1189 -5143
rect 1235 -5177 1261 -5143
rect 1303 -5177 1333 -5143
rect 1371 -5177 1405 -5143
rect 1439 -5177 1473 -5143
rect 1511 -5177 1541 -5143
rect 1583 -5177 1609 -5143
rect 1655 -5177 1677 -5143
rect 1727 -5177 1745 -5143
rect 1799 -5177 1813 -5143
rect 1871 -5177 1881 -5143
rect 1943 -5177 1949 -5143
rect 2015 -5177 2017 -5143
rect 2051 -5177 2053 -5143
rect 2119 -5177 2125 -5143
rect 2187 -5177 2197 -5143
rect 2255 -5177 2269 -5143
rect 2323 -5177 2341 -5143
rect 2391 -5177 2413 -5143
rect 2459 -5177 2485 -5143
rect 2527 -5177 2557 -5143
rect 2595 -5177 2629 -5143
rect 2663 -5177 2697 -5143
rect 2735 -5177 2790 -5143
rect -1170 -5200 2790 -5177
<< viali >>
rect -1115 -5177 -1111 -5143
rect -1111 -5177 -1081 -5143
rect -1043 -5177 -1009 -5143
rect -971 -5177 -941 -5143
rect -941 -5177 -937 -5143
rect -899 -5177 -873 -5143
rect -873 -5177 -865 -5143
rect -827 -5177 -805 -5143
rect -805 -5177 -793 -5143
rect -755 -5177 -737 -5143
rect -737 -5177 -721 -5143
rect -683 -5177 -669 -5143
rect -669 -5177 -649 -5143
rect -611 -5177 -601 -5143
rect -601 -5177 -577 -5143
rect -539 -5177 -533 -5143
rect -533 -5177 -505 -5143
rect -467 -5177 -465 -5143
rect -465 -5177 -433 -5143
rect -395 -5177 -363 -5143
rect -363 -5177 -361 -5143
rect -323 -5177 -295 -5143
rect -295 -5177 -289 -5143
rect -251 -5177 -227 -5143
rect -227 -5177 -217 -5143
rect -179 -5177 -159 -5143
rect -159 -5177 -145 -5143
rect -107 -5177 -91 -5143
rect -91 -5177 -73 -5143
rect -35 -5177 -23 -5143
rect -23 -5177 -1 -5143
rect 37 -5177 45 -5143
rect 45 -5177 71 -5143
rect 109 -5177 113 -5143
rect 113 -5177 143 -5143
rect 181 -5177 215 -5143
rect 253 -5177 283 -5143
rect 283 -5177 287 -5143
rect 325 -5177 351 -5143
rect 351 -5177 359 -5143
rect 397 -5177 419 -5143
rect 419 -5177 431 -5143
rect 469 -5177 487 -5143
rect 487 -5177 503 -5143
rect 541 -5177 555 -5143
rect 555 -5177 575 -5143
rect 613 -5177 623 -5143
rect 623 -5177 647 -5143
rect 685 -5177 691 -5143
rect 691 -5177 719 -5143
rect 757 -5177 759 -5143
rect 759 -5177 791 -5143
rect 829 -5177 861 -5143
rect 861 -5177 863 -5143
rect 901 -5177 929 -5143
rect 929 -5177 935 -5143
rect 973 -5177 997 -5143
rect 997 -5177 1007 -5143
rect 1045 -5177 1065 -5143
rect 1065 -5177 1079 -5143
rect 1117 -5177 1133 -5143
rect 1133 -5177 1151 -5143
rect 1189 -5177 1201 -5143
rect 1201 -5177 1223 -5143
rect 1261 -5177 1269 -5143
rect 1269 -5177 1295 -5143
rect 1333 -5177 1337 -5143
rect 1337 -5177 1367 -5143
rect 1405 -5177 1439 -5143
rect 1477 -5177 1507 -5143
rect 1507 -5177 1511 -5143
rect 1549 -5177 1575 -5143
rect 1575 -5177 1583 -5143
rect 1621 -5177 1643 -5143
rect 1643 -5177 1655 -5143
rect 1693 -5177 1711 -5143
rect 1711 -5177 1727 -5143
rect 1765 -5177 1779 -5143
rect 1779 -5177 1799 -5143
rect 1837 -5177 1847 -5143
rect 1847 -5177 1871 -5143
rect 1909 -5177 1915 -5143
rect 1915 -5177 1943 -5143
rect 1981 -5177 1983 -5143
rect 1983 -5177 2015 -5143
rect 2053 -5177 2085 -5143
rect 2085 -5177 2087 -5143
rect 2125 -5177 2153 -5143
rect 2153 -5177 2159 -5143
rect 2197 -5177 2221 -5143
rect 2221 -5177 2231 -5143
rect 2269 -5177 2289 -5143
rect 2289 -5177 2303 -5143
rect 2341 -5177 2357 -5143
rect 2357 -5177 2375 -5143
rect 2413 -5177 2425 -5143
rect 2425 -5177 2447 -5143
rect 2485 -5177 2493 -5143
rect 2493 -5177 2519 -5143
rect 2557 -5177 2561 -5143
rect 2561 -5177 2591 -5143
rect 2629 -5177 2663 -5143
rect 2701 -5177 2731 -5143
rect 2731 -5177 2735 -5143
<< metal1 >>
rect -1100 -3095 -780 -3080
rect -1100 -3147 -1028 -3095
rect -976 -3147 -964 -3095
rect -912 -3147 -780 -3095
rect -549 -3092 -384 -3088
rect -549 -3100 -525 -3092
rect -1100 -3160 -780 -3147
rect -580 -3144 -525 -3100
rect -473 -3144 -461 -3092
rect -409 -3100 -384 -3092
rect -53 -3094 112 -3090
rect -53 -3100 -29 -3094
rect -409 -3144 -280 -3100
rect -580 -3160 -280 -3144
rect -80 -3146 -29 -3100
rect 23 -3146 35 -3094
rect 87 -3100 112 -3094
rect 449 -3098 614 -3094
rect 1448 -3095 1613 -3091
rect 449 -3100 473 -3098
rect 87 -3146 220 -3100
rect -80 -3160 220 -3146
rect 420 -3150 473 -3100
rect 525 -3150 537 -3098
rect 589 -3100 614 -3098
rect 943 -3099 1108 -3095
rect 943 -3100 967 -3099
rect 589 -3150 720 -3100
rect 420 -3160 720 -3150
rect 920 -3151 967 -3100
rect 1019 -3151 1031 -3099
rect 1083 -3100 1108 -3099
rect 1448 -3100 1472 -3095
rect 1083 -3151 1220 -3100
rect 920 -3160 1220 -3151
rect 1420 -3147 1472 -3100
rect 1524 -3147 1536 -3095
rect 1588 -3100 1613 -3095
rect 1938 -3094 2103 -3090
rect 1588 -3147 1720 -3100
rect 1420 -3160 1720 -3147
rect 1938 -3146 1962 -3094
rect 2014 -3146 2026 -3094
rect 2078 -3100 2103 -3094
rect 2444 -3091 2609 -3087
rect 2444 -3100 2468 -3091
rect 2078 -3146 2200 -3100
rect 1938 -3150 2200 -3146
rect 1940 -3160 2200 -3150
rect 2420 -3143 2468 -3100
rect 2520 -3143 2532 -3091
rect 2584 -3100 2609 -3091
rect 2584 -3143 2720 -3100
rect 2420 -3160 2720 -3143
rect -1100 -3190 -1060 -3160
rect -1100 -3360 -1070 -3190
rect -860 -3360 -780 -3160
rect -360 -3360 -280 -3160
rect 140 -3360 220 -3160
rect 640 -3360 720 -3160
rect 1140 -3360 1220 -3160
rect 1640 -3360 1720 -3160
rect 2140 -3360 2200 -3160
rect 2640 -3360 2720 -3160
rect -1100 -3570 -780 -3360
rect -580 -3420 -280 -3360
rect -80 -3420 220 -3360
rect 420 -3420 720 -3360
rect 920 -3420 1220 -3360
rect 1420 -3420 1720 -3360
rect 1940 -3420 2200 -3360
rect 2420 -3420 2720 -3360
rect 1140 -3430 1220 -3420
rect -551 -3503 -386 -3499
rect -551 -3555 -527 -3503
rect -475 -3555 -463 -3503
rect -411 -3555 -386 -3503
rect -551 -3559 -386 -3555
rect -64 -3504 101 -3500
rect -64 -3556 -40 -3504
rect 12 -3556 24 -3504
rect 76 -3556 101 -3504
rect -64 -3560 101 -3556
rect 438 -3504 603 -3500
rect 438 -3556 462 -3504
rect 514 -3556 526 -3504
rect 578 -3556 603 -3504
rect 438 -3560 603 -3556
rect 939 -3506 1104 -3502
rect 939 -3558 963 -3506
rect 1015 -3558 1027 -3506
rect 1079 -3558 1104 -3506
rect 939 -3562 1104 -3558
rect 1448 -3504 1613 -3500
rect 1448 -3556 1472 -3504
rect 1524 -3556 1536 -3504
rect 1588 -3556 1613 -3504
rect 1448 -3560 1613 -3556
rect 1947 -3504 2112 -3500
rect 1947 -3556 1971 -3504
rect 2023 -3556 2035 -3504
rect 2087 -3556 2112 -3504
rect 1947 -3560 2112 -3556
rect 2420 -3570 2720 -3490
rect -1100 -3770 -1070 -3570
rect -860 -3770 -780 -3570
rect -350 -3644 -250 -3630
rect -350 -3696 -326 -3644
rect -274 -3696 -250 -3644
rect -350 -3710 -250 -3696
rect 150 -3644 250 -3630
rect 150 -3696 174 -3644
rect 226 -3696 250 -3644
rect 150 -3710 250 -3696
rect 650 -3644 750 -3630
rect 650 -3696 674 -3644
rect 726 -3696 750 -3644
rect 650 -3710 750 -3696
rect 1152 -3644 1240 -3629
rect 1152 -3696 1170 -3644
rect 1222 -3696 1240 -3644
rect 1152 -3710 1240 -3696
rect 1650 -3644 1750 -3630
rect 1650 -3696 1674 -3644
rect 1726 -3696 1750 -3644
rect 1650 -3710 1750 -3696
rect 2150 -3644 2250 -3630
rect 2150 -3696 2174 -3644
rect 2226 -3696 2250 -3644
rect 2150 -3710 2250 -3696
rect 2640 -3770 2720 -3570
rect -1100 -3795 -760 -3770
rect 438 -3788 603 -3784
rect -1100 -3847 -1028 -3795
rect -976 -3847 -964 -3795
rect -912 -3847 -760 -3795
rect -1100 -3870 -760 -3847
rect -564 -3795 -399 -3791
rect -564 -3847 -540 -3795
rect -488 -3847 -476 -3795
rect -424 -3847 -399 -3795
rect -564 -3851 -399 -3847
rect -57 -3792 108 -3788
rect -57 -3844 -33 -3792
rect 19 -3844 31 -3792
rect 83 -3844 108 -3792
rect 438 -3840 462 -3788
rect 514 -3840 526 -3788
rect 578 -3840 603 -3788
rect 438 -3844 603 -3840
rect 941 -3788 1106 -3784
rect 941 -3840 965 -3788
rect 1017 -3840 1029 -3788
rect 1081 -3840 1106 -3788
rect 941 -3844 1106 -3840
rect 1443 -3791 1608 -3787
rect 1443 -3843 1467 -3791
rect 1519 -3843 1531 -3791
rect 1583 -3843 1608 -3791
rect -57 -3848 108 -3844
rect 1443 -3847 1608 -3843
rect 1942 -3792 2107 -3788
rect 1942 -3844 1966 -3792
rect 2018 -3844 2030 -3792
rect 2082 -3844 2107 -3792
rect 1942 -3848 2107 -3844
rect 2420 -3795 2720 -3770
rect 2420 -3847 2469 -3795
rect 2521 -3847 2533 -3795
rect 2585 -3847 2720 -3795
rect 2420 -3850 2720 -3847
rect 2445 -3851 2610 -3850
rect -1100 -3980 -780 -3870
rect -560 -3916 -395 -3912
rect -560 -3968 -536 -3916
rect -484 -3968 -472 -3916
rect -420 -3968 -395 -3916
rect -560 -3972 -395 -3968
rect -54 -3914 111 -3910
rect 951 -3912 1116 -3908
rect -54 -3966 -30 -3914
rect 22 -3966 34 -3914
rect 86 -3966 111 -3914
rect -54 -3970 111 -3966
rect 451 -3916 616 -3912
rect 451 -3968 475 -3916
rect 527 -3968 539 -3916
rect 591 -3968 616 -3916
rect 951 -3964 975 -3912
rect 1027 -3964 1039 -3912
rect 1091 -3964 1116 -3912
rect 951 -3968 1116 -3964
rect 1445 -3915 1610 -3911
rect 1445 -3967 1472 -3915
rect 1524 -3967 1536 -3915
rect 1588 -3967 1610 -3915
rect 451 -3972 616 -3968
rect 1445 -3971 1610 -3967
rect 1947 -3912 2112 -3908
rect 1947 -3964 1971 -3912
rect 2023 -3964 2035 -3912
rect 2087 -3964 2112 -3912
rect 1947 -3968 2112 -3964
rect 2420 -3980 2720 -3900
rect -1100 -4180 -1070 -3980
rect -860 -4180 -780 -3980
rect -350 -4054 -250 -4040
rect -350 -4106 -326 -4054
rect -274 -4106 -250 -4054
rect -350 -4120 -250 -4106
rect 150 -4054 250 -4040
rect 150 -4106 174 -4054
rect 226 -4106 250 -4054
rect 150 -4120 250 -4106
rect 650 -4054 750 -4040
rect 650 -4106 674 -4054
rect 726 -4106 750 -4054
rect 650 -4120 750 -4106
rect 1150 -4054 1250 -4040
rect 1150 -4106 1174 -4054
rect 1226 -4106 1250 -4054
rect 1150 -4120 1250 -4106
rect 1650 -4054 1750 -4040
rect 1650 -4106 1674 -4054
rect 1726 -4106 1750 -4054
rect 1650 -4120 1750 -4106
rect 2150 -4054 2250 -4040
rect 2150 -4106 2174 -4054
rect 2226 -4106 2250 -4054
rect 2150 -4120 2250 -4106
rect 2640 -4180 2720 -3980
rect -1100 -4209 -780 -4180
rect -1100 -4261 -1034 -4209
rect -982 -4261 -970 -4209
rect -918 -4261 -780 -4209
rect -1100 -4390 -780 -4261
rect -556 -4208 -391 -4204
rect -556 -4260 -532 -4208
rect -480 -4260 -468 -4208
rect -416 -4260 -391 -4208
rect -556 -4264 -391 -4260
rect -55 -4205 110 -4201
rect -55 -4257 -31 -4205
rect 21 -4257 33 -4205
rect 85 -4257 110 -4205
rect -55 -4261 110 -4257
rect 445 -4204 610 -4200
rect 445 -4256 469 -4204
rect 521 -4256 533 -4204
rect 585 -4256 610 -4204
rect 1441 -4204 1606 -4200
rect 445 -4260 610 -4256
rect 937 -4215 1102 -4211
rect 937 -4267 961 -4215
rect 1013 -4267 1025 -4215
rect 1077 -4267 1102 -4215
rect 1441 -4256 1465 -4204
rect 1517 -4256 1529 -4204
rect 1581 -4256 1606 -4204
rect 1441 -4260 1606 -4256
rect 1947 -4204 2112 -4200
rect 1947 -4256 1971 -4204
rect 2023 -4256 2035 -4204
rect 2087 -4256 2112 -4204
rect 1947 -4260 2112 -4256
rect 2420 -4205 2720 -4180
rect 2420 -4257 2471 -4205
rect 2523 -4257 2535 -4205
rect 2587 -4257 2720 -4205
rect 2420 -4260 2720 -4257
rect 2447 -4261 2612 -4260
rect 937 -4271 1102 -4267
rect -552 -4323 -387 -4319
rect -552 -4375 -528 -4323
rect -476 -4375 -464 -4323
rect -412 -4375 -387 -4323
rect -552 -4379 -387 -4375
rect -61 -4325 104 -4321
rect -61 -4377 -37 -4325
rect 15 -4377 27 -4325
rect 79 -4377 104 -4325
rect -61 -4381 104 -4377
rect 453 -4323 618 -4319
rect 453 -4375 477 -4323
rect 529 -4375 541 -4323
rect 593 -4375 618 -4323
rect 453 -4379 618 -4375
rect 945 -4324 1110 -4320
rect 945 -4376 969 -4324
rect 1021 -4376 1033 -4324
rect 1085 -4376 1110 -4324
rect 945 -4380 1110 -4376
rect 1448 -4323 1613 -4319
rect 1448 -4375 1472 -4323
rect 1524 -4375 1536 -4323
rect 1588 -4375 1613 -4323
rect 1448 -4379 1613 -4375
rect 1947 -4325 2112 -4321
rect 1947 -4377 1971 -4325
rect 2023 -4377 2035 -4325
rect 2087 -4377 2112 -4325
rect 1947 -4381 2112 -4377
rect 2420 -4390 2720 -4310
rect -1100 -4590 -1070 -4390
rect -860 -4590 -780 -4390
rect -350 -4464 -250 -4450
rect -350 -4516 -326 -4464
rect -274 -4516 -250 -4464
rect -350 -4530 -250 -4516
rect 150 -4464 250 -4450
rect 150 -4516 174 -4464
rect 226 -4516 250 -4464
rect 150 -4530 250 -4516
rect 650 -4464 750 -4450
rect 650 -4516 674 -4464
rect 726 -4516 750 -4464
rect 650 -4530 750 -4516
rect 1150 -4464 1250 -4450
rect 1150 -4516 1174 -4464
rect 1226 -4516 1250 -4464
rect 1150 -4530 1250 -4516
rect 1650 -4464 1750 -4450
rect 1650 -4516 1674 -4464
rect 1726 -4516 1750 -4464
rect 1650 -4530 1750 -4516
rect 2150 -4464 2250 -4450
rect 2150 -4516 2174 -4464
rect 2226 -4516 2250 -4464
rect 2150 -4530 2250 -4516
rect 2640 -4590 2720 -4390
rect -1100 -4617 -780 -4590
rect -1100 -4669 -1034 -4617
rect -982 -4669 -970 -4617
rect -918 -4669 -780 -4617
rect -1100 -4800 -780 -4669
rect -558 -4619 -393 -4615
rect -558 -4671 -534 -4619
rect -482 -4671 -470 -4619
rect -418 -4671 -393 -4619
rect -558 -4675 -393 -4671
rect -62 -4620 103 -4616
rect -62 -4672 -38 -4620
rect 14 -4672 26 -4620
rect 78 -4672 103 -4620
rect -62 -4676 103 -4672
rect 436 -4620 601 -4616
rect 436 -4672 460 -4620
rect 512 -4672 524 -4620
rect 576 -4672 601 -4620
rect 436 -4676 601 -4672
rect 947 -4619 1112 -4615
rect 947 -4671 971 -4619
rect 1023 -4671 1035 -4619
rect 1087 -4671 1112 -4619
rect 947 -4675 1112 -4671
rect 1445 -4625 1610 -4621
rect 1445 -4677 1469 -4625
rect 1521 -4677 1533 -4625
rect 1585 -4677 1610 -4625
rect 1445 -4681 1610 -4677
rect 1938 -4624 2103 -4620
rect 1938 -4676 1962 -4624
rect 2014 -4676 2026 -4624
rect 2078 -4676 2103 -4624
rect 2420 -4623 2720 -4590
rect 2420 -4670 2467 -4623
rect 1938 -4680 2103 -4676
rect 2443 -4675 2467 -4670
rect 2519 -4675 2531 -4623
rect 2583 -4670 2720 -4623
rect 2583 -4675 2608 -4670
rect 2443 -4679 2608 -4675
rect -580 -4800 -280 -4740
rect -80 -4800 220 -4740
rect 440 -4800 720 -4740
rect 920 -4800 1220 -4740
rect 1420 -4800 1720 -4740
rect 1940 -4800 2220 -4740
rect 2420 -4800 2720 -4740
rect -1100 -5000 -1070 -4800
rect -860 -5000 -780 -4800
rect -360 -5000 -280 -4800
rect 140 -5000 220 -4800
rect 640 -5000 720 -4800
rect 1140 -5000 1220 -4800
rect 1640 -5000 1720 -4800
rect 2140 -5000 2220 -4800
rect 2640 -5000 2720 -4800
rect -1100 -5032 -780 -5000
rect -1100 -5084 -1033 -5032
rect -981 -5084 -969 -5032
rect -917 -5084 -780 -5032
rect -580 -5033 -280 -5000
rect -580 -5060 -532 -5033
rect -1100 -5120 -780 -5084
rect -556 -5085 -532 -5060
rect -480 -5085 -468 -5033
rect -416 -5060 -280 -5033
rect -80 -5028 220 -5000
rect -80 -5060 -38 -5028
rect -416 -5085 -391 -5060
rect -62 -5080 -38 -5060
rect 14 -5080 26 -5028
rect 78 -5060 220 -5028
rect 440 -5024 720 -5000
rect 440 -5060 467 -5024
rect 78 -5080 103 -5060
rect 443 -5076 467 -5060
rect 519 -5076 531 -5024
rect 583 -5060 720 -5024
rect 920 -5034 1220 -5000
rect 920 -5060 979 -5034
rect 583 -5076 608 -5060
rect 443 -5080 608 -5076
rect -62 -5084 103 -5080
rect -556 -5089 -391 -5085
rect 955 -5086 979 -5060
rect 1031 -5086 1043 -5034
rect 1095 -5060 1220 -5034
rect 1420 -5036 1720 -5000
rect 1940 -5032 2220 -5000
rect 1420 -5060 1469 -5036
rect 1095 -5086 1120 -5060
rect 955 -5090 1120 -5086
rect 1445 -5088 1469 -5060
rect 1521 -5088 1533 -5036
rect 1585 -5060 1720 -5036
rect 1937 -5036 2220 -5032
rect 1585 -5088 1610 -5060
rect 1445 -5092 1610 -5088
rect 1937 -5088 1961 -5036
rect 2013 -5088 2025 -5036
rect 2077 -5060 2220 -5036
rect 2420 -5033 2720 -5000
rect 2420 -5060 2473 -5033
rect 2077 -5088 2102 -5060
rect 1937 -5092 2102 -5088
rect 2449 -5085 2473 -5060
rect 2525 -5085 2537 -5033
rect 2589 -5060 2720 -5033
rect 2589 -5085 2614 -5060
rect 2449 -5089 2614 -5085
rect -1170 -5143 2790 -5120
rect -1170 -5177 -1115 -5143
rect -1081 -5177 -1043 -5143
rect -1009 -5177 -971 -5143
rect -937 -5177 -899 -5143
rect -865 -5177 -827 -5143
rect -793 -5177 -755 -5143
rect -721 -5177 -683 -5143
rect -649 -5177 -611 -5143
rect -577 -5177 -539 -5143
rect -505 -5177 -467 -5143
rect -433 -5177 -395 -5143
rect -361 -5177 -323 -5143
rect -289 -5177 -251 -5143
rect -217 -5177 -179 -5143
rect -145 -5177 -107 -5143
rect -73 -5177 -35 -5143
rect -1 -5177 37 -5143
rect 71 -5177 109 -5143
rect 143 -5177 181 -5143
rect 215 -5177 253 -5143
rect 287 -5177 325 -5143
rect 359 -5177 397 -5143
rect 431 -5177 469 -5143
rect 503 -5177 541 -5143
rect 575 -5177 613 -5143
rect 647 -5177 685 -5143
rect 719 -5177 757 -5143
rect 791 -5177 829 -5143
rect 863 -5177 901 -5143
rect 935 -5177 973 -5143
rect 1007 -5177 1045 -5143
rect 1079 -5177 1117 -5143
rect 1151 -5177 1189 -5143
rect 1223 -5177 1261 -5143
rect 1295 -5177 1333 -5143
rect 1367 -5177 1405 -5143
rect 1439 -5177 1477 -5143
rect 1511 -5177 1549 -5143
rect 1583 -5177 1621 -5143
rect 1655 -5177 1693 -5143
rect 1727 -5177 1765 -5143
rect 1799 -5177 1837 -5143
rect 1871 -5177 1909 -5143
rect 1943 -5177 1981 -5143
rect 2015 -5177 2053 -5143
rect 2087 -5177 2125 -5143
rect 2159 -5177 2197 -5143
rect 2231 -5177 2269 -5143
rect 2303 -5177 2341 -5143
rect 2375 -5177 2413 -5143
rect 2447 -5177 2485 -5143
rect 2519 -5177 2557 -5143
rect 2591 -5177 2629 -5143
rect 2663 -5177 2701 -5143
rect 2735 -5177 2790 -5143
rect -1170 -5200 2790 -5177
<< via1 >>
rect -1028 -3147 -976 -3095
rect -964 -3147 -912 -3095
rect -525 -3144 -473 -3092
rect -461 -3144 -409 -3092
rect -29 -3146 23 -3094
rect 35 -3146 87 -3094
rect 473 -3150 525 -3098
rect 537 -3150 589 -3098
rect 967 -3151 1019 -3099
rect 1031 -3151 1083 -3099
rect 1472 -3147 1524 -3095
rect 1536 -3147 1588 -3095
rect 1962 -3146 2014 -3094
rect 2026 -3146 2078 -3094
rect 2468 -3143 2520 -3091
rect 2532 -3143 2584 -3091
rect -527 -3555 -475 -3503
rect -463 -3555 -411 -3503
rect -40 -3556 12 -3504
rect 24 -3556 76 -3504
rect 462 -3556 514 -3504
rect 526 -3556 578 -3504
rect 963 -3558 1015 -3506
rect 1027 -3558 1079 -3506
rect 1472 -3556 1524 -3504
rect 1536 -3556 1588 -3504
rect 1971 -3556 2023 -3504
rect 2035 -3556 2087 -3504
rect -326 -3696 -274 -3644
rect 174 -3696 226 -3644
rect 674 -3696 726 -3644
rect 1170 -3696 1222 -3644
rect 1674 -3696 1726 -3644
rect 2174 -3696 2226 -3644
rect -1028 -3847 -976 -3795
rect -964 -3847 -912 -3795
rect -540 -3847 -488 -3795
rect -476 -3847 -424 -3795
rect -33 -3844 19 -3792
rect 31 -3844 83 -3792
rect 462 -3840 514 -3788
rect 526 -3840 578 -3788
rect 965 -3840 1017 -3788
rect 1029 -3840 1081 -3788
rect 1467 -3843 1519 -3791
rect 1531 -3843 1583 -3791
rect 1966 -3844 2018 -3792
rect 2030 -3844 2082 -3792
rect 2469 -3847 2521 -3795
rect 2533 -3847 2585 -3795
rect -536 -3968 -484 -3916
rect -472 -3968 -420 -3916
rect -30 -3966 22 -3914
rect 34 -3966 86 -3914
rect 475 -3968 527 -3916
rect 539 -3968 591 -3916
rect 975 -3964 1027 -3912
rect 1039 -3964 1091 -3912
rect 1472 -3967 1524 -3915
rect 1536 -3967 1588 -3915
rect 1971 -3964 2023 -3912
rect 2035 -3964 2087 -3912
rect -326 -4106 -274 -4054
rect 174 -4106 226 -4054
rect 674 -4106 726 -4054
rect 1174 -4106 1226 -4054
rect 1674 -4106 1726 -4054
rect 2174 -4106 2226 -4054
rect -1034 -4261 -982 -4209
rect -970 -4261 -918 -4209
rect -532 -4260 -480 -4208
rect -468 -4260 -416 -4208
rect -31 -4257 21 -4205
rect 33 -4257 85 -4205
rect 469 -4256 521 -4204
rect 533 -4256 585 -4204
rect 961 -4267 1013 -4215
rect 1025 -4267 1077 -4215
rect 1465 -4256 1517 -4204
rect 1529 -4256 1581 -4204
rect 1971 -4256 2023 -4204
rect 2035 -4256 2087 -4204
rect 2471 -4257 2523 -4205
rect 2535 -4257 2587 -4205
rect -528 -4375 -476 -4323
rect -464 -4375 -412 -4323
rect -37 -4377 15 -4325
rect 27 -4377 79 -4325
rect 477 -4375 529 -4323
rect 541 -4375 593 -4323
rect 969 -4376 1021 -4324
rect 1033 -4376 1085 -4324
rect 1472 -4375 1524 -4323
rect 1536 -4375 1588 -4323
rect 1971 -4377 2023 -4325
rect 2035 -4377 2087 -4325
rect -326 -4516 -274 -4464
rect 174 -4516 226 -4464
rect 674 -4516 726 -4464
rect 1174 -4516 1226 -4464
rect 1674 -4516 1726 -4464
rect 2174 -4516 2226 -4464
rect -1034 -4669 -982 -4617
rect -970 -4669 -918 -4617
rect -534 -4671 -482 -4619
rect -470 -4671 -418 -4619
rect -38 -4672 14 -4620
rect 26 -4672 78 -4620
rect 460 -4672 512 -4620
rect 524 -4672 576 -4620
rect 971 -4671 1023 -4619
rect 1035 -4671 1087 -4619
rect 1469 -4677 1521 -4625
rect 1533 -4677 1585 -4625
rect 1962 -4676 2014 -4624
rect 2026 -4676 2078 -4624
rect 2467 -4675 2519 -4623
rect 2531 -4675 2583 -4623
rect -1033 -5084 -981 -5032
rect -969 -5084 -917 -5032
rect -532 -5085 -480 -5033
rect -468 -5085 -416 -5033
rect -38 -5080 14 -5028
rect 26 -5080 78 -5028
rect 467 -5076 519 -5024
rect 531 -5076 583 -5024
rect 979 -5086 1031 -5034
rect 1043 -5086 1095 -5034
rect 1469 -5088 1521 -5036
rect 1533 -5088 1585 -5036
rect 1961 -5088 2013 -5036
rect 2025 -5088 2077 -5036
rect 2473 -5085 2525 -5033
rect 2537 -5085 2589 -5033
<< metal2 >>
rect 820 -2982 2400 -2970
rect 820 -3038 832 -2982
rect 888 -3038 2332 -2982
rect 2388 -3038 2400 -2982
rect 820 -3050 2400 -3038
rect -1060 -3091 2640 -3080
rect -1060 -3092 2468 -3091
rect -1060 -3095 -525 -3092
rect -1060 -3147 -1028 -3095
rect -976 -3147 -964 -3095
rect -912 -3144 -525 -3095
rect -473 -3144 -461 -3092
rect -409 -3094 2468 -3092
rect -409 -3144 -29 -3094
rect -912 -3146 -29 -3144
rect 23 -3146 35 -3094
rect 87 -3095 1962 -3094
rect 87 -3098 1472 -3095
rect 87 -3146 473 -3098
rect -912 -3147 473 -3146
rect -1060 -3150 473 -3147
rect 525 -3150 537 -3098
rect 589 -3099 1472 -3098
rect 589 -3150 967 -3099
rect -1060 -3151 967 -3150
rect 1019 -3151 1031 -3099
rect 1083 -3147 1472 -3099
rect 1524 -3147 1536 -3095
rect 1588 -3146 1962 -3095
rect 2014 -3146 2026 -3094
rect 2078 -3143 2468 -3094
rect 2520 -3143 2532 -3091
rect 2584 -3143 2640 -3091
rect 2078 -3146 2640 -3143
rect 1588 -3147 2640 -3146
rect 1083 -3151 2640 -3147
rect -1060 -3160 2640 -3151
rect -1042 -3161 -897 -3160
rect 459 -3164 604 -3160
rect 953 -3165 1098 -3160
rect 1458 -3161 1603 -3160
rect -541 -3490 -396 -3489
rect -172 -3490 -109 -3485
rect 827 -3490 890 -3489
rect 1829 -3490 1892 -3487
rect -580 -3501 120 -3490
rect -580 -3503 -169 -3501
rect -580 -3555 -527 -3503
rect -475 -3555 -463 -3503
rect -411 -3555 -169 -3503
rect -580 -3557 -169 -3555
rect -113 -3504 120 -3501
rect -113 -3556 -40 -3504
rect 12 -3556 24 -3504
rect 76 -3556 120 -3504
rect -113 -3557 120 -3556
rect -580 -3570 120 -3557
rect 420 -3504 1120 -3490
rect 420 -3556 462 -3504
rect 514 -3556 526 -3504
rect 578 -3505 1120 -3504
rect 578 -3556 830 -3505
rect 420 -3561 830 -3556
rect 886 -3506 1120 -3505
rect 886 -3558 963 -3506
rect 1015 -3558 1027 -3506
rect 1079 -3558 1120 -3506
rect 886 -3561 1120 -3558
rect 420 -3570 1120 -3561
rect 1420 -3503 2140 -3490
rect 1420 -3504 1832 -3503
rect 1420 -3556 1472 -3504
rect 1524 -3556 1536 -3504
rect 1588 -3556 1832 -3504
rect 1420 -3559 1832 -3556
rect 1888 -3504 2140 -3503
rect 1888 -3556 1971 -3504
rect 2023 -3556 2035 -3504
rect 2087 -3556 2140 -3504
rect 1888 -3559 2140 -3556
rect 1420 -3570 2140 -3559
rect -172 -3572 -109 -3570
rect 827 -3576 890 -3570
rect 949 -3572 1094 -3570
rect 1829 -3574 1892 -3570
rect -340 -3642 -260 -3620
rect -340 -3698 -328 -3642
rect -272 -3698 -260 -3642
rect -340 -3720 -260 -3698
rect 160 -3642 240 -3620
rect 160 -3698 172 -3642
rect 228 -3698 240 -3642
rect 160 -3720 240 -3698
rect 660 -3642 740 -3620
rect 660 -3698 672 -3642
rect 728 -3698 740 -3642
rect 660 -3720 740 -3698
rect 1162 -3642 1230 -3619
rect 1162 -3698 1168 -3642
rect 1224 -3698 1230 -3642
rect 1162 -3720 1230 -3698
rect 1660 -3642 1740 -3620
rect 1660 -3698 1672 -3642
rect 1728 -3698 1740 -3642
rect 1660 -3720 1740 -3698
rect 2160 -3642 2240 -3620
rect 2160 -3698 2172 -3642
rect 2228 -3698 2240 -3642
rect 2160 -3720 2240 -3698
rect -1042 -3790 -897 -3781
rect -554 -3790 -409 -3781
rect -47 -3790 98 -3778
rect 448 -3788 593 -3774
rect 448 -3790 462 -3788
rect -1070 -3792 462 -3790
rect -1070 -3795 -33 -3792
rect -1070 -3847 -1028 -3795
rect -976 -3847 -964 -3795
rect -912 -3847 -540 -3795
rect -488 -3847 -476 -3795
rect -424 -3844 -33 -3795
rect 19 -3844 31 -3792
rect 83 -3840 462 -3792
rect 514 -3840 526 -3788
rect 578 -3790 593 -3788
rect 951 -3788 1096 -3774
rect 951 -3790 965 -3788
rect 578 -3840 965 -3790
rect 1017 -3840 1029 -3788
rect 1081 -3790 1096 -3788
rect 1453 -3790 1598 -3777
rect 1952 -3790 2097 -3778
rect 2455 -3790 2600 -3781
rect 1081 -3791 2640 -3790
rect 1081 -3840 1467 -3791
rect 83 -3843 1467 -3840
rect 1519 -3843 1531 -3791
rect 1583 -3792 2640 -3791
rect 1583 -3843 1966 -3792
rect 83 -3844 1966 -3843
rect 2018 -3844 2030 -3792
rect 2082 -3795 2640 -3792
rect 2082 -3844 2469 -3795
rect -424 -3847 2469 -3844
rect 2521 -3847 2533 -3795
rect 2585 -3847 2640 -3795
rect -1070 -3870 2640 -3847
rect 1957 -3900 2102 -3898
rect 2312 -3900 2391 -3898
rect -580 -3912 900 -3900
rect -580 -3914 832 -3912
rect -580 -3916 -30 -3914
rect -580 -3968 -536 -3916
rect -484 -3968 -472 -3916
rect -420 -3966 -30 -3916
rect 22 -3966 34 -3914
rect 86 -3916 832 -3914
rect 86 -3966 475 -3916
rect -420 -3968 475 -3966
rect 527 -3968 539 -3916
rect 591 -3968 832 -3916
rect 888 -3968 900 -3912
rect -580 -3980 900 -3968
rect 940 -3912 1380 -3900
rect 940 -3964 975 -3912
rect 1027 -3964 1039 -3912
rect 1091 -3964 1312 -3912
rect 940 -3968 1312 -3964
rect 1368 -3968 1380 -3912
rect 940 -3980 1380 -3968
rect 1440 -3912 2400 -3900
rect 1440 -3915 1971 -3912
rect 1440 -3967 1472 -3915
rect 1524 -3967 1536 -3915
rect 1588 -3964 1971 -3915
rect 2023 -3964 2035 -3912
rect 2087 -3914 2400 -3912
rect 2087 -3964 2331 -3914
rect 1588 -3967 2331 -3964
rect 1440 -3970 2331 -3967
rect 2387 -3970 2400 -3914
rect 1440 -3980 2400 -3970
rect -550 -3982 -405 -3980
rect 461 -3982 606 -3980
rect 1455 -3981 1600 -3980
rect 2328 -3985 2391 -3980
rect -340 -4052 -260 -4030
rect -340 -4108 -328 -4052
rect -272 -4108 -260 -4052
rect -340 -4130 -260 -4108
rect 160 -4052 240 -4030
rect 160 -4108 172 -4052
rect 228 -4108 240 -4052
rect 160 -4130 240 -4108
rect 660 -4052 740 -4030
rect 660 -4108 672 -4052
rect 728 -4108 740 -4052
rect 660 -4130 740 -4108
rect 1160 -4052 1240 -4030
rect 1160 -4108 1172 -4052
rect 1228 -4108 1240 -4052
rect 1160 -4130 1240 -4108
rect 1660 -4052 1740 -4030
rect 1660 -4108 1672 -4052
rect 1728 -4108 1740 -4052
rect 1660 -4130 1740 -4108
rect 2160 -4052 2240 -4030
rect 2160 -4108 2172 -4052
rect 2228 -4108 2240 -4052
rect 2160 -4130 2240 -4108
rect -1048 -4200 -903 -4195
rect -546 -4200 -401 -4194
rect -45 -4200 100 -4191
rect 455 -4200 600 -4190
rect 1451 -4200 1596 -4190
rect 1957 -4200 2102 -4190
rect 2457 -4200 2602 -4191
rect -1080 -4204 2640 -4200
rect -1080 -4205 469 -4204
rect -1080 -4208 -31 -4205
rect -1080 -4209 -532 -4208
rect -1080 -4261 -1034 -4209
rect -982 -4261 -970 -4209
rect -918 -4260 -532 -4209
rect -480 -4260 -468 -4208
rect -416 -4257 -31 -4208
rect 21 -4257 33 -4205
rect 85 -4256 469 -4205
rect 521 -4256 533 -4204
rect 585 -4215 1465 -4204
rect 585 -4256 961 -4215
rect 85 -4257 961 -4256
rect -416 -4260 961 -4257
rect -918 -4261 961 -4260
rect -1080 -4267 961 -4261
rect 1013 -4267 1025 -4215
rect 1077 -4256 1465 -4215
rect 1517 -4256 1529 -4204
rect 1581 -4256 1971 -4204
rect 2023 -4256 2035 -4204
rect 2087 -4205 2640 -4204
rect 2087 -4256 2471 -4205
rect 1077 -4257 2471 -4256
rect 2523 -4257 2535 -4205
rect 2587 -4257 2640 -4205
rect 1077 -4267 2640 -4257
rect -1080 -4280 2640 -4267
rect -542 -4310 -397 -4309
rect -170 -4310 -107 -4308
rect 463 -4310 608 -4309
rect 1458 -4310 1603 -4309
rect -580 -4323 120 -4310
rect -580 -4375 -528 -4323
rect -476 -4375 -464 -4323
rect -412 -4324 120 -4323
rect -412 -4375 -167 -4324
rect -580 -4380 -167 -4375
rect -111 -4325 120 -4324
rect -111 -4377 -37 -4325
rect 15 -4377 27 -4325
rect 79 -4377 120 -4325
rect -111 -4380 120 -4377
rect -580 -4390 120 -4380
rect 420 -4322 1140 -4310
rect 420 -4323 832 -4322
rect 420 -4375 477 -4323
rect 529 -4375 541 -4323
rect 593 -4375 832 -4323
rect 420 -4378 832 -4375
rect 888 -4324 1140 -4322
rect 888 -4376 969 -4324
rect 1021 -4376 1033 -4324
rect 1085 -4376 1140 -4324
rect 888 -4378 1140 -4376
rect 420 -4390 1140 -4378
rect 1420 -4322 2120 -4310
rect 1420 -4323 1832 -4322
rect 1420 -4375 1472 -4323
rect 1524 -4375 1536 -4323
rect 1588 -4375 1832 -4323
rect 1420 -4378 1832 -4375
rect 1888 -4325 2120 -4322
rect 1888 -4377 1971 -4325
rect 2023 -4377 2035 -4325
rect 2087 -4377 2120 -4325
rect 1888 -4378 2120 -4377
rect 1420 -4390 2120 -4378
rect -170 -4395 -107 -4390
rect -51 -4391 94 -4390
rect 1957 -4391 2102 -4390
rect -340 -4462 -260 -4440
rect -340 -4518 -328 -4462
rect -272 -4518 -260 -4462
rect -340 -4540 -260 -4518
rect 160 -4462 240 -4440
rect 160 -4518 172 -4462
rect 228 -4518 240 -4462
rect 160 -4540 240 -4518
rect 660 -4462 740 -4440
rect 660 -4518 672 -4462
rect 728 -4518 740 -4462
rect 660 -4540 740 -4518
rect 1160 -4462 1240 -4440
rect 1160 -4518 1172 -4462
rect 1228 -4518 1240 -4462
rect 1160 -4540 1240 -4518
rect 1660 -4462 1740 -4440
rect 1660 -4518 1672 -4462
rect 1728 -4518 1740 -4462
rect 1660 -4540 1740 -4518
rect 2160 -4462 2240 -4440
rect 2160 -4518 2172 -4462
rect 2228 -4518 2240 -4462
rect 2160 -4540 2240 -4518
rect -1048 -4610 -903 -4603
rect -548 -4610 -403 -4605
rect -52 -4610 93 -4606
rect 446 -4610 591 -4606
rect 957 -4610 1102 -4605
rect 2453 -4610 2598 -4609
rect -1070 -4617 2640 -4610
rect -1070 -4669 -1034 -4617
rect -982 -4669 -970 -4617
rect -918 -4619 2640 -4617
rect -918 -4669 -534 -4619
rect -1070 -4671 -534 -4669
rect -482 -4671 -470 -4619
rect -418 -4620 971 -4619
rect -418 -4671 -38 -4620
rect -1070 -4672 -38 -4671
rect 14 -4672 26 -4620
rect 78 -4672 460 -4620
rect 512 -4672 524 -4620
rect 576 -4671 971 -4620
rect 1023 -4671 1035 -4619
rect 1087 -4623 2640 -4619
rect 1087 -4624 2467 -4623
rect 1087 -4625 1962 -4624
rect 1087 -4671 1469 -4625
rect 576 -4672 1469 -4671
rect -1070 -4677 1469 -4672
rect 1521 -4677 1533 -4625
rect 1585 -4676 1962 -4625
rect 2014 -4676 2026 -4624
rect 2078 -4675 2467 -4624
rect 2519 -4675 2531 -4623
rect 2583 -4675 2640 -4623
rect 2078 -4676 2640 -4675
rect 1585 -4677 2640 -4676
rect -1070 -4690 2640 -4677
rect -1047 -5020 -902 -5018
rect -546 -5020 -401 -5019
rect -52 -5020 93 -5014
rect 453 -5020 598 -5010
rect 2459 -5020 2604 -5019
rect -1070 -5024 2640 -5020
rect -1070 -5028 467 -5024
rect -1070 -5032 -38 -5028
rect -1070 -5084 -1033 -5032
rect -981 -5084 -969 -5032
rect -917 -5033 -38 -5032
rect -917 -5084 -532 -5033
rect -1070 -5085 -532 -5084
rect -480 -5085 -468 -5033
rect -416 -5080 -38 -5033
rect 14 -5080 26 -5028
rect 78 -5076 467 -5028
rect 519 -5076 531 -5024
rect 583 -5033 2640 -5024
rect 583 -5034 2473 -5033
rect 583 -5076 979 -5034
rect 78 -5080 979 -5076
rect -416 -5085 979 -5080
rect -1070 -5086 979 -5085
rect 1031 -5086 1043 -5034
rect 1095 -5036 2473 -5034
rect 1095 -5086 1469 -5036
rect -1070 -5088 1469 -5086
rect 1521 -5088 1533 -5036
rect 1585 -5088 1961 -5036
rect 2013 -5088 2025 -5036
rect 2077 -5085 2473 -5036
rect 2525 -5085 2537 -5033
rect 2589 -5085 2640 -5033
rect 2077 -5088 2640 -5085
rect -1070 -5100 2640 -5088
rect 1455 -5102 1600 -5100
rect 1947 -5102 2092 -5100
<< via2 >>
rect 832 -3038 888 -2982
rect 2332 -3038 2388 -2982
rect -169 -3557 -113 -3501
rect 830 -3561 886 -3505
rect 1832 -3559 1888 -3503
rect -328 -3644 -272 -3642
rect -328 -3696 -326 -3644
rect -326 -3696 -274 -3644
rect -274 -3696 -272 -3644
rect -328 -3698 -272 -3696
rect 172 -3644 228 -3642
rect 172 -3696 174 -3644
rect 174 -3696 226 -3644
rect 226 -3696 228 -3644
rect 172 -3698 228 -3696
rect 672 -3644 728 -3642
rect 672 -3696 674 -3644
rect 674 -3696 726 -3644
rect 726 -3696 728 -3644
rect 672 -3698 728 -3696
rect 1168 -3644 1224 -3642
rect 1168 -3696 1170 -3644
rect 1170 -3696 1222 -3644
rect 1222 -3696 1224 -3644
rect 1168 -3698 1224 -3696
rect 1672 -3644 1728 -3642
rect 1672 -3696 1674 -3644
rect 1674 -3696 1726 -3644
rect 1726 -3696 1728 -3644
rect 1672 -3698 1728 -3696
rect 2172 -3644 2228 -3642
rect 2172 -3696 2174 -3644
rect 2174 -3696 2226 -3644
rect 2226 -3696 2228 -3644
rect 2172 -3698 2228 -3696
rect 832 -3968 888 -3912
rect 1312 -3968 1368 -3912
rect 2331 -3970 2387 -3914
rect -328 -4054 -272 -4052
rect -328 -4106 -326 -4054
rect -326 -4106 -274 -4054
rect -274 -4106 -272 -4054
rect -328 -4108 -272 -4106
rect 172 -4054 228 -4052
rect 172 -4106 174 -4054
rect 174 -4106 226 -4054
rect 226 -4106 228 -4054
rect 172 -4108 228 -4106
rect 672 -4054 728 -4052
rect 672 -4106 674 -4054
rect 674 -4106 726 -4054
rect 726 -4106 728 -4054
rect 672 -4108 728 -4106
rect 1172 -4054 1228 -4052
rect 1172 -4106 1174 -4054
rect 1174 -4106 1226 -4054
rect 1226 -4106 1228 -4054
rect 1172 -4108 1228 -4106
rect 1672 -4054 1728 -4052
rect 1672 -4106 1674 -4054
rect 1674 -4106 1726 -4054
rect 1726 -4106 1728 -4054
rect 1672 -4108 1728 -4106
rect 2172 -4054 2228 -4052
rect 2172 -4106 2174 -4054
rect 2174 -4106 2226 -4054
rect 2226 -4106 2228 -4054
rect 2172 -4108 2228 -4106
rect -167 -4380 -111 -4324
rect 832 -4378 888 -4322
rect 1832 -4378 1888 -4322
rect -328 -4464 -272 -4462
rect -328 -4516 -326 -4464
rect -326 -4516 -274 -4464
rect -274 -4516 -272 -4464
rect -328 -4518 -272 -4516
rect 172 -4464 228 -4462
rect 172 -4516 174 -4464
rect 174 -4516 226 -4464
rect 226 -4516 228 -4464
rect 172 -4518 228 -4516
rect 672 -4464 728 -4462
rect 672 -4516 674 -4464
rect 674 -4516 726 -4464
rect 726 -4516 728 -4464
rect 672 -4518 728 -4516
rect 1172 -4464 1228 -4462
rect 1172 -4516 1174 -4464
rect 1174 -4516 1226 -4464
rect 1226 -4516 1228 -4464
rect 1172 -4518 1228 -4516
rect 1672 -4464 1728 -4462
rect 1672 -4516 1674 -4464
rect 1674 -4516 1726 -4464
rect 1726 -4516 1728 -4464
rect 1672 -4518 1728 -4516
rect 2172 -4464 2228 -4462
rect 2172 -4516 2174 -4464
rect 2174 -4516 2226 -4464
rect 2226 -4516 2228 -4464
rect 2172 -4518 2228 -4516
<< metal3 >>
rect 820 -2982 900 -2970
rect 820 -3038 832 -2982
rect 888 -3038 900 -2982
rect -180 -3423 -90 -3410
rect -180 -3487 -167 -3423
rect -103 -3487 -90 -3423
rect -180 -3490 -90 -3487
rect -182 -3500 -90 -3490
rect 820 -3494 900 -3038
rect 1800 -3070 1900 -2890
rect 1820 -3410 1900 -3070
rect 2320 -2982 2400 -2890
rect 2320 -3038 2332 -2982
rect 2388 -3038 2400 -2982
rect -182 -3501 -99 -3500
rect -182 -3557 -169 -3501
rect -113 -3557 -99 -3501
rect -182 -3567 -99 -3557
rect 817 -3505 900 -3494
rect 817 -3561 830 -3505
rect 886 -3561 900 -3505
rect -340 -3625 -260 -3590
rect -350 -3638 -250 -3625
rect -350 -3702 -332 -3638
rect -268 -3702 -250 -3638
rect -350 -3715 -250 -3702
rect -340 -3750 -260 -3715
rect -340 -4035 -260 -4020
rect -350 -4048 -250 -4035
rect -350 -4112 -332 -4048
rect -268 -4112 -250 -4048
rect -350 -4125 -250 -4112
rect -340 -4160 -260 -4125
rect -180 -4313 -100 -3567
rect 817 -3571 900 -3561
rect 160 -3625 240 -3590
rect 660 -3625 740 -3590
rect 150 -3638 250 -3625
rect 150 -3702 168 -3638
rect 232 -3702 250 -3638
rect 150 -3715 250 -3702
rect 650 -3638 750 -3625
rect 650 -3702 668 -3638
rect 732 -3702 750 -3638
rect 650 -3715 750 -3702
rect 160 -3750 240 -3715
rect 660 -3750 740 -3715
rect 820 -3899 900 -3571
rect 1300 -3423 1390 -3410
rect 1300 -3487 1313 -3423
rect 1377 -3487 1390 -3423
rect 1300 -3500 1390 -3487
rect 1820 -3423 1910 -3410
rect 1820 -3487 1828 -3423
rect 1892 -3487 1910 -3423
rect 1820 -3492 1910 -3487
rect 1819 -3500 1910 -3492
rect 1140 -3638 1240 -3590
rect 1140 -3702 1158 -3638
rect 1222 -3642 1240 -3638
rect 1224 -3698 1240 -3642
rect 1222 -3702 1240 -3698
rect 1140 -3750 1240 -3702
rect 818 -3912 901 -3899
rect 818 -3968 832 -3912
rect 888 -3968 901 -3912
rect 818 -3976 901 -3968
rect 1300 -3912 1380 -3500
rect 1819 -3503 1902 -3500
rect 1819 -3559 1832 -3503
rect 1888 -3559 1902 -3503
rect 1819 -3569 1902 -3559
rect 1660 -3625 1740 -3590
rect 1650 -3638 1750 -3625
rect 1650 -3702 1668 -3638
rect 1732 -3702 1750 -3638
rect 1650 -3715 1750 -3702
rect 1660 -3750 1740 -3715
rect 1300 -3968 1312 -3912
rect 1368 -3968 1380 -3912
rect 160 -4035 240 -4020
rect 660 -4035 740 -4020
rect 150 -4048 250 -4035
rect 150 -4112 168 -4048
rect 232 -4112 250 -4048
rect 150 -4125 250 -4112
rect 650 -4048 750 -4035
rect 650 -4112 668 -4048
rect 732 -4112 750 -4048
rect 650 -4125 750 -4112
rect 160 -4160 240 -4125
rect 660 -4160 740 -4125
rect -180 -4324 -97 -4313
rect -180 -4380 -167 -4324
rect -111 -4380 -97 -4324
rect -180 -4390 -97 -4380
rect 820 -4322 900 -3976
rect 1300 -3980 1380 -3968
rect 1160 -4035 1240 -4020
rect 1660 -4035 1740 -4020
rect 1150 -4048 1250 -4035
rect 1150 -4112 1168 -4048
rect 1232 -4112 1250 -4048
rect 1150 -4125 1250 -4112
rect 1650 -4048 1750 -4035
rect 1650 -4112 1668 -4048
rect 1732 -4112 1750 -4048
rect 1650 -4125 1750 -4112
rect 1160 -4160 1240 -4125
rect 1660 -4160 1740 -4125
rect 820 -4378 832 -4322
rect 888 -4378 900 -4322
rect 820 -4390 900 -4378
rect 1820 -4322 1900 -3569
rect 2160 -3625 2240 -3590
rect 2150 -3638 2250 -3625
rect 2150 -3702 2168 -3638
rect 2232 -3702 2250 -3638
rect 2150 -3715 2250 -3702
rect 2160 -3750 2240 -3715
rect 2320 -3903 2400 -3038
rect 2640 -3643 2720 -3630
rect 2640 -3707 2653 -3643
rect 2717 -3707 2720 -3643
rect 2318 -3914 2401 -3903
rect 2318 -3970 2331 -3914
rect 2387 -3970 2401 -3914
rect 2318 -3980 2401 -3970
rect 2160 -4035 2240 -4020
rect 2640 -4030 2720 -3707
rect 2150 -4048 2250 -4035
rect 2150 -4112 2168 -4048
rect 2232 -4112 2250 -4048
rect 2150 -4125 2250 -4112
rect 2640 -4043 2730 -4030
rect 2640 -4107 2653 -4043
rect 2717 -4107 2730 -4043
rect 2640 -4120 2730 -4107
rect 2160 -4160 2240 -4125
rect 1820 -4378 1832 -4322
rect 1888 -4378 1900 -4322
rect 1820 -4390 1900 -4378
rect -340 -4445 -260 -4430
rect 160 -4445 240 -4410
rect 660 -4445 740 -4430
rect 1160 -4445 1240 -4430
rect 1660 -4445 1740 -4430
rect 2160 -4445 2240 -4430
rect 2640 -4440 2720 -4120
rect -350 -4458 -250 -4445
rect -350 -4522 -332 -4458
rect -268 -4522 -250 -4458
rect -350 -4535 -250 -4522
rect 150 -4458 250 -4445
rect 150 -4522 168 -4458
rect 232 -4522 250 -4458
rect 150 -4535 250 -4522
rect 650 -4458 750 -4445
rect 650 -4522 668 -4458
rect 732 -4522 750 -4458
rect 650 -4535 750 -4522
rect 1150 -4458 1250 -4445
rect 1150 -4522 1168 -4458
rect 1232 -4522 1250 -4458
rect 1150 -4535 1250 -4522
rect 1650 -4458 1750 -4445
rect 1650 -4522 1668 -4458
rect 1732 -4522 1750 -4458
rect 1650 -4535 1750 -4522
rect 2150 -4458 2250 -4445
rect 2150 -4522 2168 -4458
rect 2232 -4522 2250 -4458
rect 2150 -4535 2250 -4522
rect 2640 -4453 2730 -4440
rect 2640 -4517 2653 -4453
rect 2717 -4517 2730 -4453
rect 2640 -4530 2730 -4517
rect -340 -4570 -260 -4535
rect 160 -4570 240 -4535
rect 660 -4570 740 -4535
rect 1160 -4570 1240 -4535
rect 1660 -4570 1740 -4535
rect 2160 -4570 2240 -4535
<< via3 >>
rect -167 -3487 -103 -3423
rect -332 -3642 -268 -3638
rect -332 -3698 -328 -3642
rect -328 -3698 -272 -3642
rect -272 -3698 -268 -3642
rect -332 -3702 -268 -3698
rect -332 -4052 -268 -4048
rect -332 -4108 -328 -4052
rect -328 -4108 -272 -4052
rect -272 -4108 -268 -4052
rect -332 -4112 -268 -4108
rect 168 -3642 232 -3638
rect 168 -3698 172 -3642
rect 172 -3698 228 -3642
rect 228 -3698 232 -3642
rect 168 -3702 232 -3698
rect 668 -3642 732 -3638
rect 668 -3698 672 -3642
rect 672 -3698 728 -3642
rect 728 -3698 732 -3642
rect 668 -3702 732 -3698
rect 1313 -3487 1377 -3423
rect 1828 -3487 1892 -3423
rect 1158 -3642 1222 -3638
rect 1158 -3698 1168 -3642
rect 1168 -3698 1222 -3642
rect 1158 -3702 1222 -3698
rect 1668 -3642 1732 -3638
rect 1668 -3698 1672 -3642
rect 1672 -3698 1728 -3642
rect 1728 -3698 1732 -3642
rect 1668 -3702 1732 -3698
rect 168 -4052 232 -4048
rect 168 -4108 172 -4052
rect 172 -4108 228 -4052
rect 228 -4108 232 -4052
rect 168 -4112 232 -4108
rect 668 -4052 732 -4048
rect 668 -4108 672 -4052
rect 672 -4108 728 -4052
rect 728 -4108 732 -4052
rect 668 -4112 732 -4108
rect 1168 -4052 1232 -4048
rect 1168 -4108 1172 -4052
rect 1172 -4108 1228 -4052
rect 1228 -4108 1232 -4052
rect 1168 -4112 1232 -4108
rect 1668 -4052 1732 -4048
rect 1668 -4108 1672 -4052
rect 1672 -4108 1728 -4052
rect 1728 -4108 1732 -4052
rect 1668 -4112 1732 -4108
rect 2168 -3642 2232 -3638
rect 2168 -3698 2172 -3642
rect 2172 -3698 2228 -3642
rect 2228 -3698 2232 -3642
rect 2168 -3702 2232 -3698
rect 2653 -3707 2717 -3643
rect 2168 -4052 2232 -4048
rect 2168 -4108 2172 -4052
rect 2172 -4108 2228 -4052
rect 2228 -4108 2232 -4052
rect 2168 -4112 2232 -4108
rect 2653 -4107 2717 -4043
rect -332 -4462 -268 -4458
rect -332 -4518 -328 -4462
rect -328 -4518 -272 -4462
rect -272 -4518 -268 -4462
rect -332 -4522 -268 -4518
rect 168 -4462 232 -4458
rect 168 -4518 172 -4462
rect 172 -4518 228 -4462
rect 228 -4518 232 -4462
rect 168 -4522 232 -4518
rect 668 -4462 732 -4458
rect 668 -4518 672 -4462
rect 672 -4518 728 -4462
rect 728 -4518 732 -4462
rect 668 -4522 732 -4518
rect 1168 -4462 1232 -4458
rect 1168 -4518 1172 -4462
rect 1172 -4518 1228 -4462
rect 1228 -4518 1232 -4462
rect 1168 -4522 1232 -4518
rect 1668 -4462 1732 -4458
rect 1668 -4518 1672 -4462
rect 1672 -4518 1728 -4462
rect 1728 -4518 1732 -4462
rect 1668 -4522 1732 -4518
rect 2168 -4462 2232 -4458
rect 2168 -4518 2172 -4462
rect 2172 -4518 2228 -4462
rect 2228 -4518 2232 -4462
rect 2168 -4522 2232 -4518
rect 2653 -4517 2717 -4453
<< metal4 >>
rect -180 -3423 1910 -3410
rect -180 -3487 -167 -3423
rect -103 -3487 1313 -3423
rect 1377 -3487 1828 -3423
rect 1892 -3487 1910 -3423
rect -180 -3500 1910 -3487
rect -341 -3630 -259 -3629
rect 159 -3630 241 -3629
rect 659 -3630 741 -3629
rect 1149 -3630 1231 -3629
rect 1659 -3630 1741 -3629
rect 2159 -3630 2241 -3629
rect -1070 -3638 2790 -3630
rect -1070 -3702 -332 -3638
rect -268 -3702 168 -3638
rect 232 -3702 668 -3638
rect 732 -3702 1158 -3638
rect 1222 -3702 1668 -3638
rect 1732 -3702 2168 -3638
rect 2232 -3643 2790 -3638
rect 2232 -3702 2653 -3643
rect -1070 -3707 2653 -3702
rect 2717 -3707 2790 -3643
rect -1070 -3710 2790 -3707
rect -341 -3711 -259 -3710
rect 159 -3711 241 -3710
rect 659 -3711 741 -3710
rect 1149 -3711 1231 -3710
rect 1659 -3711 1741 -3710
rect 2159 -3711 2241 -3710
rect 2640 -3720 2790 -3710
rect -341 -4040 -259 -4039
rect 159 -4040 241 -4039
rect 659 -4040 741 -4039
rect 1159 -4040 1241 -4039
rect 1659 -4040 1741 -4039
rect 2159 -4040 2241 -4039
rect 2640 -4040 2730 -4030
rect -1070 -4043 2730 -4040
rect -1070 -4048 2653 -4043
rect -1070 -4112 -332 -4048
rect -268 -4112 168 -4048
rect 232 -4112 668 -4048
rect 732 -4112 1168 -4048
rect 1232 -4112 1668 -4048
rect 1732 -4112 2168 -4048
rect 2232 -4107 2653 -4048
rect 2717 -4107 2730 -4043
rect 2232 -4112 2730 -4107
rect -1070 -4120 2730 -4112
rect -341 -4121 -259 -4120
rect 159 -4121 241 -4120
rect 659 -4121 741 -4120
rect 1159 -4121 1241 -4120
rect 1659 -4121 1741 -4120
rect 2159 -4121 2241 -4120
rect 2640 -4121 2720 -4120
rect -341 -4450 -259 -4449
rect 159 -4450 241 -4449
rect 659 -4450 741 -4449
rect 1159 -4450 1241 -4449
rect 1659 -4450 1741 -4449
rect 2159 -4450 2241 -4449
rect 2640 -4450 2730 -4440
rect -1070 -4453 2730 -4450
rect -1070 -4458 2653 -4453
rect -1070 -4522 -332 -4458
rect -268 -4522 168 -4458
rect 232 -4522 668 -4458
rect 732 -4522 1168 -4458
rect 1232 -4522 1668 -4458
rect 1732 -4522 2168 -4458
rect 2232 -4517 2653 -4458
rect 2717 -4517 2730 -4453
rect 2232 -4522 2730 -4517
rect -1070 -4530 2730 -4522
rect -341 -4531 -259 -4530
rect 159 -4531 241 -4530
rect 659 -4531 741 -4530
rect 1159 -4531 1241 -4530
rect 1659 -4531 1741 -4530
rect 2159 -4531 2241 -4530
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_0
timestamp 1757161594
transform 0 1 57 -1 0 -3672
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_1
timestamp 1757161594
transform 0 1 -943 -1 0 -3262
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_2
timestamp 1757161594
transform 0 1 -443 -1 0 -3262
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_3
timestamp 1757161594
transform 0 1 57 -1 0 -3262
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_4
timestamp 1757161594
transform 0 1 557 -1 0 -3262
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_5
timestamp 1757161594
transform 0 1 1057 -1 0 -3262
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_6
timestamp 1757161594
transform 0 1 1557 -1 0 -3262
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_7
timestamp 1757161594
transform 0 1 2057 -1 0 -3262
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_8
timestamp 1757161594
transform 0 1 2557 -1 0 -3262
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_9
timestamp 1757161594
transform 0 1 -943 -1 0 -3672
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_10
timestamp 1757161594
transform 0 1 -443 -1 0 -3672
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_11
timestamp 1757161594
transform 0 1 1057 -1 0 -3672
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_12
timestamp 1757161594
transform 0 1 557 -1 0 -3672
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_13
timestamp 1757161594
transform 0 1 2057 -1 0 -3672
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_14
timestamp 1757161594
transform 0 1 1557 -1 0 -3672
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_15
timestamp 1757161594
transform 0 1 57 -1 0 -4082
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_16
timestamp 1757161594
transform 0 1 2557 -1 0 -3672
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_17
timestamp 1757161594
transform 0 1 -943 -1 0 -4082
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_18
timestamp 1757161594
transform 0 1 -443 -1 0 -4082
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_19
timestamp 1757161594
transform 0 1 1057 -1 0 -4082
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_20
timestamp 1757161594
transform 0 1 557 -1 0 -4082
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_21
timestamp 1757161594
transform 0 1 2057 -1 0 -4082
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_22
timestamp 1757161594
transform 0 1 1557 -1 0 -4082
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_23
timestamp 1757161594
transform 0 1 57 -1 0 -4492
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_24
timestamp 1757161594
transform 0 1 2557 -1 0 -4082
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_25
timestamp 1757161594
transform 0 1 -943 -1 0 -4492
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_26
timestamp 1757161594
transform 0 1 -443 -1 0 -4492
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_27
timestamp 1757161594
transform 0 1 1057 -1 0 -4492
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_28
timestamp 1757161594
transform 0 1 557 -1 0 -4492
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_29
timestamp 1757161594
transform 0 1 2057 -1 0 -4492
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_30
timestamp 1757161594
transform 0 1 1557 -1 0 -4492
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_31
timestamp 1757161594
transform 0 1 57 -1 0 -4902
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_32
timestamp 1757161594
transform 0 1 2557 -1 0 -4492
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_33
timestamp 1757161594
transform 0 1 -943 -1 0 -4902
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_34
timestamp 1757161594
transform 0 1 -443 -1 0 -4902
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_35
timestamp 1757161594
transform 0 1 1057 -1 0 -4902
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_36
timestamp 1757161594
transform 0 1 557 -1 0 -4902
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_37
timestamp 1757161594
transform 0 1 2057 -1 0 -4902
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_38
timestamp 1757161594
transform 0 1 1557 -1 0 -4902
box -184 -157 184 157
use sky130_fd_pr__nfet_01v8_lvt_34DASA  sky130_fd_pr__nfet_01v8_lvt_34DASA_39
timestamp 1757161594
transform 0 1 2557 -1 0 -4902
box -184 -157 184 157
<< end >>
