magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -194 -298 194 264
<< pmoslvt >>
rect -100 -236 100 164
<< pdiff >>
rect -158 151 -100 164
rect -158 117 -146 151
rect -112 117 -100 151
rect -158 83 -100 117
rect -158 49 -146 83
rect -112 49 -100 83
rect -158 15 -100 49
rect -158 -19 -146 15
rect -112 -19 -100 15
rect -158 -53 -100 -19
rect -158 -87 -146 -53
rect -112 -87 -100 -53
rect -158 -121 -100 -87
rect -158 -155 -146 -121
rect -112 -155 -100 -121
rect -158 -189 -100 -155
rect -158 -223 -146 -189
rect -112 -223 -100 -189
rect -158 -236 -100 -223
rect 100 151 158 164
rect 100 117 112 151
rect 146 117 158 151
rect 100 83 158 117
rect 100 49 112 83
rect 146 49 158 83
rect 100 15 158 49
rect 100 -19 112 15
rect 146 -19 158 15
rect 100 -53 158 -19
rect 100 -87 112 -53
rect 146 -87 158 -53
rect 100 -121 158 -87
rect 100 -155 112 -121
rect 146 -155 158 -121
rect 100 -189 158 -155
rect 100 -223 112 -189
rect 146 -223 158 -189
rect 100 -236 158 -223
<< pdiffc >>
rect -146 117 -112 151
rect -146 49 -112 83
rect -146 -19 -112 15
rect -146 -87 -112 -53
rect -146 -155 -112 -121
rect -146 -223 -112 -189
rect 112 117 146 151
rect 112 49 146 83
rect 112 -19 146 15
rect 112 -87 146 -53
rect 112 -155 146 -121
rect 112 -223 146 -189
<< poly >>
rect -100 245 100 261
rect -100 211 -51 245
rect -17 211 17 245
rect 51 211 100 245
rect -100 164 100 211
rect -100 -262 100 -236
<< polycont >>
rect -51 211 -17 245
rect 17 211 51 245
<< locali >>
rect -100 211 -53 245
rect -17 211 17 245
rect 53 211 100 245
rect -146 151 -112 168
rect -146 83 -112 91
rect -146 15 -112 19
rect -146 -91 -112 -87
rect -146 -163 -112 -155
rect -146 -240 -112 -223
rect 112 151 146 168
rect 112 83 146 91
rect 112 15 146 19
rect 112 -91 146 -87
rect 112 -163 146 -155
rect 112 -240 146 -223
<< viali >>
rect -53 211 -51 245
rect -51 211 -19 245
rect 19 211 51 245
rect 51 211 53 245
rect -146 117 -112 125
rect -146 91 -112 117
rect -146 49 -112 53
rect -146 19 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -91
rect -146 -125 -112 -121
rect -146 -189 -112 -163
rect -146 -197 -112 -189
rect 112 117 146 125
rect 112 91 146 117
rect 112 49 146 53
rect 112 19 146 49
rect 112 -53 146 -19
rect 112 -121 146 -91
rect 112 -125 146 -121
rect 112 -189 146 -163
rect 112 -197 146 -189
<< metal1 >>
rect -96 245 96 251
rect -96 211 -53 245
rect -19 211 19 245
rect 53 211 96 245
rect -96 205 96 211
rect -152 125 -106 164
rect -152 91 -146 125
rect -112 91 -106 125
rect -152 53 -106 91
rect -152 19 -146 53
rect -112 19 -106 53
rect -152 -19 -106 19
rect -152 -53 -146 -19
rect -112 -53 -106 -19
rect -152 -91 -106 -53
rect -152 -125 -146 -91
rect -112 -125 -106 -91
rect -152 -163 -106 -125
rect -152 -197 -146 -163
rect -112 -197 -106 -163
rect -152 -236 -106 -197
rect 106 125 152 164
rect 106 91 112 125
rect 146 91 152 125
rect 106 53 152 91
rect 106 19 112 53
rect 146 19 152 53
rect 106 -19 152 19
rect 106 -53 112 -19
rect 146 -53 152 -19
rect 106 -91 152 -53
rect 106 -125 112 -91
rect 146 -125 152 -91
rect 106 -163 152 -125
rect 106 -197 112 -163
rect 146 -197 152 -163
rect 106 -236 152 -197
<< end >>
