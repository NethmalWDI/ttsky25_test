magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< metal3 >>
rect -686 992 686 1040
rect -686 928 602 992
rect 666 928 686 992
rect -686 912 686 928
rect -686 848 602 912
rect 666 848 686 912
rect -686 832 686 848
rect -686 768 602 832
rect 666 768 686 832
rect -686 752 686 768
rect -686 688 602 752
rect 666 688 686 752
rect -686 672 686 688
rect -686 608 602 672
rect 666 608 686 672
rect -686 592 686 608
rect -686 528 602 592
rect 666 528 686 592
rect -686 512 686 528
rect -686 448 602 512
rect 666 448 686 512
rect -686 432 686 448
rect -686 368 602 432
rect 666 368 686 432
rect -686 352 686 368
rect -686 288 602 352
rect 666 288 686 352
rect -686 272 686 288
rect -686 208 602 272
rect 666 208 686 272
rect -686 192 686 208
rect -686 128 602 192
rect 666 128 686 192
rect -686 112 686 128
rect -686 48 602 112
rect 666 48 686 112
rect -686 32 686 48
rect -686 -32 602 32
rect 666 -32 686 32
rect -686 -48 686 -32
rect -686 -112 602 -48
rect 666 -112 686 -48
rect -686 -128 686 -112
rect -686 -192 602 -128
rect 666 -192 686 -128
rect -686 -208 686 -192
rect -686 -272 602 -208
rect 666 -272 686 -208
rect -686 -288 686 -272
rect -686 -352 602 -288
rect 666 -352 686 -288
rect -686 -368 686 -352
rect -686 -432 602 -368
rect 666 -432 686 -368
rect -686 -448 686 -432
rect -686 -512 602 -448
rect 666 -512 686 -448
rect -686 -528 686 -512
rect -686 -592 602 -528
rect 666 -592 686 -528
rect -686 -608 686 -592
rect -686 -672 602 -608
rect 666 -672 686 -608
rect -686 -688 686 -672
rect -686 -752 602 -688
rect 666 -752 686 -688
rect -686 -768 686 -752
rect -686 -832 602 -768
rect 666 -832 686 -768
rect -686 -848 686 -832
rect -686 -912 602 -848
rect 666 -912 686 -848
rect -686 -928 686 -912
rect -686 -992 602 -928
rect 666 -992 686 -928
rect -686 -1040 686 -992
<< via3 >>
rect 602 928 666 992
rect 602 848 666 912
rect 602 768 666 832
rect 602 688 666 752
rect 602 608 666 672
rect 602 528 666 592
rect 602 448 666 512
rect 602 368 666 432
rect 602 288 666 352
rect 602 208 666 272
rect 602 128 666 192
rect 602 48 666 112
rect 602 -32 666 32
rect 602 -112 666 -48
rect 602 -192 666 -128
rect 602 -272 666 -208
rect 602 -352 666 -288
rect 602 -432 666 -368
rect 602 -512 666 -448
rect 602 -592 666 -528
rect 602 -672 666 -608
rect 602 -752 666 -688
rect 602 -832 666 -768
rect 602 -912 666 -848
rect 602 -992 666 -928
<< mimcap >>
rect -646 952 354 1000
rect -646 -952 -578 952
rect 286 -952 354 952
rect -646 -1000 354 -952
<< mimcapcontact >>
rect -578 -952 286 952
<< metal4 >>
rect 586 992 682 1028
rect -607 952 315 961
rect -607 -952 -578 952
rect 286 -952 315 952
rect -607 -961 315 -952
rect 586 928 602 992
rect 666 928 682 992
rect 586 912 682 928
rect 586 848 602 912
rect 666 848 682 912
rect 586 832 682 848
rect 586 768 602 832
rect 666 768 682 832
rect 586 752 682 768
rect 586 688 602 752
rect 666 688 682 752
rect 586 672 682 688
rect 586 608 602 672
rect 666 608 682 672
rect 586 592 682 608
rect 586 528 602 592
rect 666 528 682 592
rect 586 512 682 528
rect 586 448 602 512
rect 666 448 682 512
rect 586 432 682 448
rect 586 368 602 432
rect 666 368 682 432
rect 586 352 682 368
rect 586 288 602 352
rect 666 288 682 352
rect 586 272 682 288
rect 586 208 602 272
rect 666 208 682 272
rect 586 192 682 208
rect 586 128 602 192
rect 666 128 682 192
rect 586 112 682 128
rect 586 48 602 112
rect 666 48 682 112
rect 586 32 682 48
rect 586 -32 602 32
rect 666 -32 682 32
rect 586 -48 682 -32
rect 586 -112 602 -48
rect 666 -112 682 -48
rect 586 -128 682 -112
rect 586 -192 602 -128
rect 666 -192 682 -128
rect 586 -208 682 -192
rect 586 -272 602 -208
rect 666 -272 682 -208
rect 586 -288 682 -272
rect 586 -352 602 -288
rect 666 -352 682 -288
rect 586 -368 682 -352
rect 586 -432 602 -368
rect 666 -432 682 -368
rect 586 -448 682 -432
rect 586 -512 602 -448
rect 666 -512 682 -448
rect 586 -528 682 -512
rect 586 -592 602 -528
rect 666 -592 682 -528
rect 586 -608 682 -592
rect 586 -672 602 -608
rect 666 -672 682 -608
rect 586 -688 682 -672
rect 586 -752 602 -688
rect 666 -752 682 -688
rect 586 -768 682 -752
rect 586 -832 602 -768
rect 666 -832 682 -768
rect 586 -848 682 -832
rect 586 -912 602 -848
rect 666 -912 682 -848
rect 586 -928 682 -912
rect 586 -992 602 -928
rect 666 -992 682 -928
rect 586 -1028 682 -992
<< properties >>
string FIXED_BBOX -686 -1040 394 1040
<< end >>
