magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -1094 -148 1094 114
<< pmoslvt >>
rect -1000 -86 1000 14
<< pdiff >>
rect -1058 -19 -1000 14
rect -1058 -53 -1046 -19
rect -1012 -53 -1000 -19
rect -1058 -86 -1000 -53
rect 1000 -19 1058 14
rect 1000 -53 1012 -19
rect 1046 -53 1058 -19
rect 1000 -86 1058 -53
<< pdiffc >>
rect -1046 -53 -1012 -19
rect 1012 -53 1046 -19
<< poly >>
rect -705 95 705 111
rect -705 78 -663 95
rect -1000 61 -663 78
rect -629 61 -595 95
rect -561 61 -527 95
rect -493 61 -459 95
rect -425 61 -391 95
rect -357 61 -323 95
rect -289 61 -255 95
rect -221 61 -187 95
rect -153 61 -119 95
rect -85 61 -51 95
rect -17 61 17 95
rect 51 61 85 95
rect 119 61 153 95
rect 187 61 221 95
rect 255 61 289 95
rect 323 61 357 95
rect 391 61 425 95
rect 459 61 493 95
rect 527 61 561 95
rect 595 61 629 95
rect 663 78 705 95
rect 663 61 1000 78
rect -1000 14 1000 61
rect -1000 -112 1000 -86
<< polycont >>
rect -663 61 -629 95
rect -595 61 -561 95
rect -527 61 -493 95
rect -459 61 -425 95
rect -391 61 -357 95
rect -323 61 -289 95
rect -255 61 -221 95
rect -187 61 -153 95
rect -119 61 -85 95
rect -51 61 -17 95
rect 17 61 51 95
rect 85 61 119 95
rect 153 61 187 95
rect 221 61 255 95
rect 289 61 323 95
rect 357 61 391 95
rect 425 61 459 95
rect 493 61 527 95
rect 561 61 595 95
rect 629 61 663 95
<< locali >>
rect -705 61 -665 95
rect -629 61 -595 95
rect -559 61 -527 95
rect -487 61 -459 95
rect -415 61 -391 95
rect -343 61 -323 95
rect -271 61 -255 95
rect -199 61 -187 95
rect -127 61 -119 95
rect -55 61 -51 95
rect 51 61 55 95
rect 119 61 127 95
rect 187 61 199 95
rect 255 61 271 95
rect 323 61 343 95
rect 391 61 415 95
rect 459 61 487 95
rect 527 61 559 95
rect 595 61 629 95
rect 665 61 705 95
rect -1046 -19 -1012 7
rect -1046 -79 -1012 -53
rect 1012 -19 1046 7
rect 1012 -79 1046 -53
<< viali >>
rect -665 61 -663 95
rect -663 61 -631 95
rect -593 61 -561 95
rect -561 61 -559 95
rect -521 61 -493 95
rect -493 61 -487 95
rect -449 61 -425 95
rect -425 61 -415 95
rect -377 61 -357 95
rect -357 61 -343 95
rect -305 61 -289 95
rect -289 61 -271 95
rect -233 61 -221 95
rect -221 61 -199 95
rect -161 61 -153 95
rect -153 61 -127 95
rect -89 61 -85 95
rect -85 61 -55 95
rect -17 61 17 95
rect 55 61 85 95
rect 85 61 89 95
rect 127 61 153 95
rect 153 61 161 95
rect 199 61 221 95
rect 221 61 233 95
rect 271 61 289 95
rect 289 61 305 95
rect 343 61 357 95
rect 357 61 377 95
rect 415 61 425 95
rect 425 61 449 95
rect 487 61 493 95
rect 493 61 521 95
rect 559 61 561 95
rect 561 61 593 95
rect 631 61 663 95
rect 663 61 665 95
rect -1046 -53 -1012 -19
rect 1012 -53 1046 -19
<< metal1 >>
rect -701 95 701 101
rect -701 61 -665 95
rect -631 61 -593 95
rect -559 61 -521 95
rect -487 61 -449 95
rect -415 61 -377 95
rect -343 61 -305 95
rect -271 61 -233 95
rect -199 61 -161 95
rect -127 61 -89 95
rect -55 61 -17 95
rect 17 61 55 95
rect 89 61 127 95
rect 161 61 199 95
rect 233 61 271 95
rect 305 61 343 95
rect 377 61 415 95
rect 449 61 487 95
rect 521 61 559 95
rect 593 61 631 95
rect 665 61 701 95
rect -701 55 701 61
rect -1052 -19 -1006 3
rect -1052 -53 -1046 -19
rect -1012 -53 -1006 -19
rect -1052 -75 -1006 -53
rect 1006 -19 1052 3
rect 1006 -53 1012 -19
rect 1046 -53 1052 -19
rect 1006 -75 1052 -53
<< end >>
