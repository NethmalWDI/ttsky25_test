magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -286 -369 286 369
<< nmoslvt >>
rect -100 -169 100 231
<< ndiff >>
rect -158 218 -100 231
rect -158 184 -146 218
rect -112 184 -100 218
rect -158 150 -100 184
rect -158 116 -146 150
rect -112 116 -100 150
rect -158 82 -100 116
rect -158 48 -146 82
rect -112 48 -100 82
rect -158 14 -100 48
rect -158 -20 -146 14
rect -112 -20 -100 14
rect -158 -54 -100 -20
rect -158 -88 -146 -54
rect -112 -88 -100 -54
rect -158 -122 -100 -88
rect -158 -156 -146 -122
rect -112 -156 -100 -122
rect -158 -169 -100 -156
rect 100 218 158 231
rect 100 184 112 218
rect 146 184 158 218
rect 100 150 158 184
rect 100 116 112 150
rect 146 116 158 150
rect 100 82 158 116
rect 100 48 112 82
rect 146 48 158 82
rect 100 14 158 48
rect 100 -20 112 14
rect 146 -20 158 14
rect 100 -54 158 -20
rect 100 -88 112 -54
rect 146 -88 158 -54
rect 100 -122 158 -88
rect 100 -156 112 -122
rect 146 -156 158 -122
rect 100 -169 158 -156
<< ndiffc >>
rect -146 184 -112 218
rect -146 116 -112 150
rect -146 48 -112 82
rect -146 -20 -112 14
rect -146 -88 -112 -54
rect -146 -156 -112 -122
rect 112 184 146 218
rect 112 116 146 150
rect 112 48 146 82
rect 112 -20 146 14
rect 112 -88 146 -54
rect 112 -156 146 -122
<< psubdiff >>
rect -260 309 260 343
rect -260 -309 -226 309
rect 226 221 260 309
rect 226 153 260 187
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect 226 -119 260 -85
rect 226 -187 260 -153
rect 226 -309 260 -221
rect -260 -343 260 -309
<< psubdiffcont >>
rect 226 187 260 221
rect 226 119 260 153
rect 226 51 260 85
rect 226 -17 260 17
rect 226 -85 260 -51
rect 226 -153 260 -119
rect 226 -221 260 -187
<< poly >>
rect -100 231 100 257
rect -100 -207 100 -169
rect -100 -241 -51 -207
rect -17 -241 17 -207
rect 51 -241 100 -207
rect -100 -257 100 -241
<< polycont >>
rect -51 -241 -17 -207
rect 17 -241 51 -207
<< locali >>
rect -260 309 260 343
rect -260 -309 -226 309
rect -146 218 -112 235
rect -146 150 -112 158
rect -146 82 -112 86
rect -146 -24 -112 -20
rect -146 -96 -112 -88
rect -146 -173 -112 -156
rect 112 218 146 235
rect 112 150 146 158
rect 112 82 146 86
rect 112 -24 146 -20
rect 112 -96 146 -88
rect 112 -173 146 -156
rect 226 221 260 309
rect 226 153 260 187
rect 226 85 260 119
rect 226 17 260 51
rect 226 -51 260 -17
rect 226 -119 260 -85
rect 226 -187 260 -153
rect -100 -241 -53 -207
rect -17 -241 17 -207
rect 53 -241 100 -207
rect 226 -309 260 -221
rect -260 -343 260 -309
<< viali >>
rect -146 184 -112 192
rect -146 158 -112 184
rect -146 116 -112 120
rect -146 86 -112 116
rect -146 14 -112 48
rect -146 -54 -112 -24
rect -146 -58 -112 -54
rect -146 -122 -112 -96
rect -146 -130 -112 -122
rect 112 184 146 192
rect 112 158 146 184
rect 112 116 146 120
rect 112 86 146 116
rect 112 14 146 48
rect 112 -54 146 -24
rect 112 -58 146 -54
rect 112 -122 146 -96
rect 112 -130 146 -122
rect -53 -241 -51 -207
rect -51 -241 -19 -207
rect 19 -241 51 -207
rect 51 -241 53 -207
<< metal1 >>
rect -152 192 -106 231
rect -152 158 -146 192
rect -112 158 -106 192
rect -152 120 -106 158
rect -152 86 -146 120
rect -112 86 -106 120
rect -152 48 -106 86
rect -152 14 -146 48
rect -112 14 -106 48
rect -152 -24 -106 14
rect -152 -58 -146 -24
rect -112 -58 -106 -24
rect -152 -96 -106 -58
rect -152 -130 -146 -96
rect -112 -130 -106 -96
rect -152 -169 -106 -130
rect 106 192 152 231
rect 106 158 112 192
rect 146 158 152 192
rect 106 120 152 158
rect 106 86 112 120
rect 146 86 152 120
rect 106 48 152 86
rect 106 14 112 48
rect 146 14 152 48
rect 106 -24 152 14
rect 106 -58 112 -24
rect 146 -58 152 -24
rect 106 -96 152 -58
rect 106 -130 112 -96
rect 146 -130 152 -96
rect 106 -169 152 -130
rect -96 -207 96 -201
rect -96 -241 -53 -207
rect -19 -241 19 -207
rect 53 -241 96 -207
rect -96 -247 96 -241
<< properties >>
string FIXED_BBOX -243 -326 243 326
<< end >>
