magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< error_s >>
rect 12420 23083 12450 23181
rect 12166 23047 12565 23083
rect 12326 23013 12397 23047
rect 12363 23011 12397 23013
rect 12364 22607 12397 23011
rect 12400 23013 12588 23047
rect 12400 22977 12486 23013
rect 12400 22643 12433 22977
rect 12880 18867 13064 19004
rect 12790 18750 12810 18838
rect 12890 18750 13064 18867
rect 12810 18670 13064 18750
rect 12226 18110 12440 18364
rect 12442 18030 12670 18198
rect 12890 18030 12924 18364
rect 12480 17590 12648 18030
rect 12226 17280 12440 17534
rect 12480 17280 12610 17348
rect 12670 17280 12800 17348
rect 12480 17180 12648 17280
rect 12670 17180 12838 17280
rect 12890 17180 13054 17534
rect 12364 16393 12397 16396
rect 12400 16357 12433 16360
rect 22690 13830 22730 13891
rect 22690 13770 22790 13811
rect -6570 987 -6500 1020
rect -6570 923 -6567 987
rect -6510 923 -6500 987
rect -6570 890 -6500 923
rect -6450 987 -6380 1020
rect -6450 923 -6440 987
rect -6450 890 -6380 923
<< nwell >>
rect 5390 21830 5740 21850
rect 5390 21500 5400 21830
rect 5720 21500 5740 21830
rect 12790 18670 12810 18750
rect 17450 18280 17900 18880
rect 17450 18230 17920 18280
rect 12480 18030 12670 18110
rect 12480 17590 12610 18030
rect 12480 17180 12610 17280
rect 12670 17180 12800 17280
rect -610 16180 -570 16660
rect 17630 16350 17920 18230
<< pwell >>
rect 20244 14454 20356 14556
rect 20674 14453 20786 14456
rect 20674 14367 22113 14453
rect 20674 14364 20786 14367
rect 8647 12927 10623 13013
rect 8647 11613 8733 12927
rect 10537 11613 10623 12927
rect 20674 12676 20766 14364
rect 20674 12673 20786 12676
rect 22027 12673 22113 14367
rect 20674 12587 22113 12673
rect 20674 12584 20786 12587
rect 8647 11527 10623 11613
<< psubdiff >>
rect 20270 14480 20330 14530
rect 20700 14427 20760 14430
rect 20700 14393 20805 14427
rect 20839 14393 20873 14427
rect 20907 14393 20941 14427
rect 20975 14393 21009 14427
rect 21043 14393 21077 14427
rect 21111 14393 21145 14427
rect 21179 14393 21213 14427
rect 21247 14393 21281 14427
rect 21315 14393 21349 14427
rect 21383 14393 21417 14427
rect 21451 14393 21485 14427
rect 21519 14393 21553 14427
rect 21587 14393 21621 14427
rect 21655 14393 21689 14427
rect 21723 14393 21757 14427
rect 21791 14393 21825 14427
rect 21859 14393 21893 14427
rect 21927 14393 21961 14427
rect 21995 14393 22087 14427
rect 20700 14390 20760 14393
rect 8673 12953 8734 12987
rect 8768 12953 8802 12987
rect 8836 12953 8870 12987
rect 8904 12953 8938 12987
rect 8972 12953 9006 12987
rect 9040 12953 9074 12987
rect 9108 12953 9142 12987
rect 9176 12953 9210 12987
rect 9244 12953 9278 12987
rect 9312 12953 9346 12987
rect 9380 12953 9414 12987
rect 9448 12953 9482 12987
rect 9516 12953 9550 12987
rect 9584 12953 9618 12987
rect 9652 12953 9686 12987
rect 9720 12953 9754 12987
rect 9788 12953 9822 12987
rect 9856 12953 9890 12987
rect 9924 12953 9958 12987
rect 9992 12953 10026 12987
rect 10060 12953 10094 12987
rect 10128 12953 10162 12987
rect 10196 12953 10230 12987
rect 10264 12953 10298 12987
rect 10332 12953 10366 12987
rect 10400 12953 10434 12987
rect 10468 12953 10502 12987
rect 10536 12953 10597 12987
rect 8673 12899 8707 12953
rect 8673 12831 8707 12865
rect 8673 12763 8707 12797
rect 8673 12695 8707 12729
rect 8673 12627 8707 12661
rect 8673 12559 8707 12593
rect 8673 12491 8707 12525
rect 8673 12423 8707 12457
rect 8673 12355 8707 12389
rect 8673 12287 8707 12321
rect 8673 12219 8707 12253
rect 8673 12151 8707 12185
rect 8673 12083 8707 12117
rect 8673 12015 8707 12049
rect 8673 11947 8707 11981
rect 8673 11879 8707 11913
rect 8673 11811 8707 11845
rect 8673 11743 8707 11777
rect 8673 11675 8707 11709
rect 8673 11587 8707 11641
rect 10563 12899 10597 12953
rect 10563 12831 10597 12865
rect 10563 12763 10597 12797
rect 10563 12695 10597 12729
rect 10563 12627 10597 12661
rect 20700 12650 20740 14390
rect 22053 14353 22087 14393
rect 22053 14285 22087 14319
rect 22053 14217 22087 14251
rect 22053 14149 22087 14183
rect 22053 14081 22087 14115
rect 22053 14013 22087 14047
rect 22053 13945 22087 13979
rect 22053 13877 22087 13911
rect 22053 13809 22087 13843
rect 22053 13741 22087 13775
rect 22053 13673 22087 13707
rect 22053 13605 22087 13639
rect 22053 13537 22087 13571
rect 22053 13469 22087 13503
rect 22053 13401 22087 13435
rect 22053 13333 22087 13367
rect 22053 13265 22087 13299
rect 22053 13197 22087 13231
rect 22053 13129 22087 13163
rect 22053 13061 22087 13095
rect 22053 12993 22087 13027
rect 22053 12925 22087 12959
rect 22053 12857 22087 12891
rect 22053 12789 22087 12823
rect 22053 12721 22087 12755
rect 20700 12647 20760 12650
rect 22053 12647 22087 12687
rect 20700 12613 20805 12647
rect 20839 12613 20873 12647
rect 20907 12613 20941 12647
rect 20975 12613 21009 12647
rect 21043 12613 21077 12647
rect 21111 12613 21145 12647
rect 21179 12613 21213 12647
rect 21247 12613 21281 12647
rect 21315 12613 21349 12647
rect 21383 12613 21417 12647
rect 21451 12613 21485 12647
rect 21519 12613 21553 12647
rect 21587 12613 21621 12647
rect 21655 12613 21689 12647
rect 21723 12613 21757 12647
rect 21791 12613 21825 12647
rect 21859 12613 21893 12647
rect 21927 12613 21961 12647
rect 21995 12613 22087 12647
rect 20700 12610 20760 12613
rect 10563 12559 10597 12593
rect 10563 12491 10597 12525
rect 10563 12423 10597 12457
rect 10563 12355 10597 12389
rect 10563 12287 10597 12321
rect 10563 12219 10597 12253
rect 10563 12151 10597 12185
rect 10563 12083 10597 12117
rect 10563 12015 10597 12049
rect 10563 11947 10597 11981
rect 10563 11879 10597 11913
rect 10563 11811 10597 11845
rect 10563 11743 10597 11777
rect 10563 11675 10597 11709
rect 10563 11587 10597 11641
rect 8673 11553 8734 11587
rect 8768 11553 8802 11587
rect 8836 11553 8870 11587
rect 8904 11553 8938 11587
rect 8972 11553 9006 11587
rect 9040 11553 9074 11587
rect 9108 11553 9142 11587
rect 9176 11553 9210 11587
rect 9244 11553 9278 11587
rect 9312 11553 9346 11587
rect 9380 11553 9414 11587
rect 9448 11553 9482 11587
rect 9516 11553 9550 11587
rect 9584 11553 9618 11587
rect 9652 11553 9686 11587
rect 9720 11553 9754 11587
rect 9788 11553 9822 11587
rect 9856 11553 9890 11587
rect 9924 11553 9958 11587
rect 9992 11553 10026 11587
rect 10060 11553 10094 11587
rect 10128 11553 10162 11587
rect 10196 11553 10230 11587
rect 10264 11553 10298 11587
rect 10332 11553 10366 11587
rect 10400 11553 10434 11587
rect 10468 11553 10502 11587
rect 10536 11553 10597 11587
<< psubdiffcont >>
rect 20805 14393 20839 14427
rect 20873 14393 20907 14427
rect 20941 14393 20975 14427
rect 21009 14393 21043 14427
rect 21077 14393 21111 14427
rect 21145 14393 21179 14427
rect 21213 14393 21247 14427
rect 21281 14393 21315 14427
rect 21349 14393 21383 14427
rect 21417 14393 21451 14427
rect 21485 14393 21519 14427
rect 21553 14393 21587 14427
rect 21621 14393 21655 14427
rect 21689 14393 21723 14427
rect 21757 14393 21791 14427
rect 21825 14393 21859 14427
rect 21893 14393 21927 14427
rect 21961 14393 21995 14427
rect 8734 12953 8768 12987
rect 8802 12953 8836 12987
rect 8870 12953 8904 12987
rect 8938 12953 8972 12987
rect 9006 12953 9040 12987
rect 9074 12953 9108 12987
rect 9142 12953 9176 12987
rect 9210 12953 9244 12987
rect 9278 12953 9312 12987
rect 9346 12953 9380 12987
rect 9414 12953 9448 12987
rect 9482 12953 9516 12987
rect 9550 12953 9584 12987
rect 9618 12953 9652 12987
rect 9686 12953 9720 12987
rect 9754 12953 9788 12987
rect 9822 12953 9856 12987
rect 9890 12953 9924 12987
rect 9958 12953 9992 12987
rect 10026 12953 10060 12987
rect 10094 12953 10128 12987
rect 10162 12953 10196 12987
rect 10230 12953 10264 12987
rect 10298 12953 10332 12987
rect 10366 12953 10400 12987
rect 10434 12953 10468 12987
rect 10502 12953 10536 12987
rect 8673 12865 8707 12899
rect 8673 12797 8707 12831
rect 8673 12729 8707 12763
rect 8673 12661 8707 12695
rect 8673 12593 8707 12627
rect 8673 12525 8707 12559
rect 8673 12457 8707 12491
rect 8673 12389 8707 12423
rect 8673 12321 8707 12355
rect 8673 12253 8707 12287
rect 8673 12185 8707 12219
rect 8673 12117 8707 12151
rect 8673 12049 8707 12083
rect 8673 11981 8707 12015
rect 8673 11913 8707 11947
rect 8673 11845 8707 11879
rect 8673 11777 8707 11811
rect 8673 11709 8707 11743
rect 8673 11641 8707 11675
rect 10563 12865 10597 12899
rect 10563 12797 10597 12831
rect 10563 12729 10597 12763
rect 10563 12661 10597 12695
rect 10563 12593 10597 12627
rect 22053 14319 22087 14353
rect 22053 14251 22087 14285
rect 22053 14183 22087 14217
rect 22053 14115 22087 14149
rect 22053 14047 22087 14081
rect 22053 13979 22087 14013
rect 22053 13911 22087 13945
rect 22053 13843 22087 13877
rect 22053 13775 22087 13809
rect 22053 13707 22087 13741
rect 22053 13639 22087 13673
rect 22053 13571 22087 13605
rect 22053 13503 22087 13537
rect 22053 13435 22087 13469
rect 22053 13367 22087 13401
rect 22053 13299 22087 13333
rect 22053 13231 22087 13265
rect 22053 13163 22087 13197
rect 22053 13095 22087 13129
rect 22053 13027 22087 13061
rect 22053 12959 22087 12993
rect 22053 12891 22087 12925
rect 22053 12823 22087 12857
rect 22053 12755 22087 12789
rect 22053 12687 22087 12721
rect 20805 12613 20839 12647
rect 20873 12613 20907 12647
rect 20941 12613 20975 12647
rect 21009 12613 21043 12647
rect 21077 12613 21111 12647
rect 21145 12613 21179 12647
rect 21213 12613 21247 12647
rect 21281 12613 21315 12647
rect 21349 12613 21383 12647
rect 21417 12613 21451 12647
rect 21485 12613 21519 12647
rect 21553 12613 21587 12647
rect 21621 12613 21655 12647
rect 21689 12613 21723 12647
rect 21757 12613 21791 12647
rect 21825 12613 21859 12647
rect 21893 12613 21927 12647
rect 21961 12613 21995 12647
rect 10563 12525 10597 12559
rect 10563 12457 10597 12491
rect 10563 12389 10597 12423
rect 10563 12321 10597 12355
rect 10563 12253 10597 12287
rect 10563 12185 10597 12219
rect 10563 12117 10597 12151
rect 10563 12049 10597 12083
rect 10563 11981 10597 12015
rect 10563 11913 10597 11947
rect 10563 11845 10597 11879
rect 10563 11777 10597 11811
rect 10563 11709 10597 11743
rect 10563 11641 10597 11675
rect 8734 11553 8768 11587
rect 8802 11553 8836 11587
rect 8870 11553 8904 11587
rect 8938 11553 8972 11587
rect 9006 11553 9040 11587
rect 9074 11553 9108 11587
rect 9142 11553 9176 11587
rect 9210 11553 9244 11587
rect 9278 11553 9312 11587
rect 9346 11553 9380 11587
rect 9414 11553 9448 11587
rect 9482 11553 9516 11587
rect 9550 11553 9584 11587
rect 9618 11553 9652 11587
rect 9686 11553 9720 11587
rect 9754 11553 9788 11587
rect 9822 11553 9856 11587
rect 9890 11553 9924 11587
rect 9958 11553 9992 11587
rect 10026 11553 10060 11587
rect 10094 11553 10128 11587
rect 10162 11553 10196 11587
rect 10230 11553 10264 11587
rect 10298 11553 10332 11587
rect 10366 11553 10400 11587
rect 10434 11553 10468 11587
rect 10502 11553 10536 11587
<< locali >>
rect 20270 14480 20330 14530
rect 20700 14427 20760 14430
rect 20700 14393 20805 14427
rect 20839 14393 20873 14427
rect 20907 14393 20941 14427
rect 20975 14393 21009 14427
rect 21043 14393 21077 14427
rect 21111 14393 21145 14427
rect 21179 14393 21213 14427
rect 21247 14393 21281 14427
rect 21315 14393 21349 14427
rect 21383 14393 21417 14427
rect 21451 14393 21485 14427
rect 21519 14393 21553 14427
rect 21587 14393 21621 14427
rect 21655 14393 21689 14427
rect 21723 14393 21757 14427
rect 21791 14393 21825 14427
rect 21859 14393 21893 14427
rect 21927 14393 21961 14427
rect 21995 14393 22087 14427
rect 20700 14390 20760 14393
rect 8673 12953 8734 12987
rect 8768 12953 8802 12987
rect 8836 12953 8870 12987
rect 8904 12953 8938 12987
rect 8972 12953 9006 12987
rect 9040 12953 9074 12987
rect 9108 12953 9142 12987
rect 9176 12953 9210 12987
rect 9244 12953 9278 12987
rect 9312 12953 9346 12987
rect 9380 12953 9414 12987
rect 9448 12953 9482 12987
rect 9516 12953 9550 12987
rect 9584 12953 9618 12987
rect 9652 12953 9686 12987
rect 9720 12953 9754 12987
rect 9788 12953 9822 12987
rect 9856 12953 9890 12987
rect 9924 12953 9958 12987
rect 9992 12953 10026 12987
rect 10060 12953 10094 12987
rect 10128 12953 10162 12987
rect 10196 12953 10230 12987
rect 10264 12953 10298 12987
rect 10332 12953 10366 12987
rect 10400 12953 10434 12987
rect 10468 12953 10502 12987
rect 10536 12953 10597 12987
rect 8673 12899 8707 12953
rect 8673 12831 8707 12865
rect 8673 12763 8707 12797
rect 8673 12695 8707 12729
rect 8673 12627 8707 12661
rect 8673 12559 8707 12593
rect 8673 12491 8707 12525
rect 8673 12423 8707 12457
rect 8673 12355 8707 12389
rect 8673 12287 8707 12321
rect 8673 12219 8707 12253
rect 8673 12151 8707 12185
rect 8673 12083 8707 12117
rect 8673 12015 8707 12049
rect 8673 11947 8707 11981
rect 8673 11879 8707 11913
rect 8673 11811 8707 11845
rect 8673 11743 8707 11777
rect 8673 11675 8707 11709
rect 8673 11587 8707 11641
rect 10563 12899 10597 12953
rect 10563 12831 10597 12865
rect 10563 12763 10597 12797
rect 10563 12695 10597 12729
rect 10563 12627 10597 12661
rect 20700 12650 20740 14390
rect 22053 14353 22087 14393
rect 22053 14285 22087 14319
rect 22053 14217 22087 14251
rect 22053 14149 22087 14183
rect 22053 14081 22087 14115
rect 22053 14013 22087 14047
rect 22053 13945 22087 13979
rect 22053 13877 22087 13911
rect 22053 13809 22087 13843
rect 22053 13741 22087 13775
rect 22053 13673 22087 13707
rect 22053 13605 22087 13639
rect 22053 13537 22087 13571
rect 22053 13469 22087 13503
rect 22053 13401 22087 13435
rect 22053 13333 22087 13367
rect 22053 13265 22087 13299
rect 22053 13197 22087 13231
rect 22053 13129 22087 13163
rect 22053 13061 22087 13095
rect 22053 12993 22087 13027
rect 22053 12925 22087 12959
rect 22053 12857 22087 12891
rect 22053 12789 22087 12823
rect 22053 12721 22087 12755
rect 20700 12647 20760 12650
rect 22053 12647 22087 12687
rect 20700 12613 20805 12647
rect 20839 12613 20873 12647
rect 20907 12613 20941 12647
rect 20975 12613 21009 12647
rect 21043 12613 21077 12647
rect 21111 12613 21145 12647
rect 21179 12613 21213 12647
rect 21247 12613 21281 12647
rect 21315 12613 21349 12647
rect 21383 12613 21417 12647
rect 21451 12613 21485 12647
rect 21519 12613 21553 12647
rect 21587 12613 21621 12647
rect 21655 12613 21689 12647
rect 21723 12613 21757 12647
rect 21791 12613 21825 12647
rect 21859 12613 21893 12647
rect 21927 12613 21961 12647
rect 21995 12613 22087 12647
rect 20700 12610 20760 12613
rect 10563 12559 10597 12593
rect 10563 12491 10597 12525
rect 10563 12423 10597 12457
rect 10563 12355 10597 12389
rect 10563 12287 10597 12321
rect 10563 12219 10597 12253
rect 10563 12151 10597 12185
rect 10563 12083 10597 12117
rect 10563 12015 10597 12049
rect 10563 11947 10597 11981
rect 10563 11879 10597 11913
rect 10563 11811 10597 11845
rect 10563 11743 10597 11777
rect 10563 11675 10597 11709
rect 10563 11587 10597 11641
rect 8673 11553 8734 11587
rect 8768 11553 8802 11587
rect 8836 11553 8870 11587
rect 8904 11553 8938 11587
rect 8972 11553 9006 11587
rect 9040 11553 9074 11587
rect 9108 11553 9142 11587
rect 9176 11553 9210 11587
rect 9244 11553 9278 11587
rect 9312 11553 9346 11587
rect 9380 11553 9414 11587
rect 9448 11553 9482 11587
rect 9516 11553 9550 11587
rect 9584 11553 9618 11587
rect 9652 11553 9686 11587
rect 9720 11553 9754 11587
rect 9788 11553 9822 11587
rect 9856 11553 9890 11587
rect 9924 11553 9958 11587
rect 9992 11553 10026 11587
rect 10060 11553 10094 11587
rect 10128 11553 10162 11587
rect 10196 11553 10230 11587
rect 10264 11553 10298 11587
rect 10332 11553 10366 11587
rect 10400 11553 10434 11587
rect 10468 11553 10502 11587
rect 10536 11553 10597 11587
<< metal1 >>
rect -10440 25266 -10080 25300
rect -10440 25214 -10411 25266
rect -10359 25214 -10286 25266
rect -10234 25214 -10161 25266
rect -10109 25214 -10080 25266
rect -10440 24540 -10080 25214
rect -8670 25276 -8310 25310
rect -8670 25224 -8641 25276
rect -8589 25224 -8516 25276
rect -8464 25224 -8391 25276
rect -8339 25224 -8310 25276
rect -8670 24620 -8310 25224
rect -6940 25266 -6580 25300
rect -6940 25214 -6911 25266
rect -6859 25214 -6786 25266
rect -6734 25214 -6661 25266
rect -6609 25214 -6580 25266
rect -6940 24620 -6580 25214
rect -500 24640 -380 24650
rect -1020 24621 -380 24640
rect -1020 24569 -466 24621
rect -414 24569 -380 24621
rect -1020 24496 -380 24569
rect -1020 24444 -466 24496
rect -414 24444 -380 24496
rect -1020 24371 -380 24444
rect -1020 24340 -466 24371
rect -500 24319 -466 24340
rect -414 24319 -380 24371
rect -500 24290 -380 24319
rect -520 23431 -400 23460
rect -520 23400 -486 23431
rect -840 23379 -486 23400
rect -434 23400 -400 23431
rect -434 23379 -390 23400
rect -840 23306 -390 23379
rect -840 23254 -486 23306
rect -434 23254 -390 23306
rect -840 23181 -390 23254
rect -840 23129 -486 23181
rect -434 23129 -390 23181
rect 940 23266 1300 23300
rect 940 23214 969 23266
rect 1021 23214 1094 23266
rect 1146 23214 1219 23266
rect 1271 23214 1300 23266
rect 940 23180 1300 23214
rect 1810 23276 2170 23310
rect 1810 23224 1839 23276
rect 1891 23224 1964 23276
rect 2016 23224 2089 23276
rect 2141 23224 2170 23276
rect 1810 23190 2170 23224
rect 2710 23276 3070 23310
rect 2710 23224 2739 23276
rect 2791 23224 2864 23276
rect 2916 23224 2989 23276
rect 3041 23224 3070 23276
rect 2710 23190 3070 23224
rect 3610 23276 3970 23310
rect 3610 23224 3639 23276
rect 3691 23224 3764 23276
rect 3816 23224 3889 23276
rect 3941 23224 3970 23276
rect 3610 23190 3970 23224
rect 4500 23276 4860 23310
rect 4500 23224 4529 23276
rect 4581 23224 4654 23276
rect 4706 23224 4779 23276
rect 4831 23224 4860 23276
rect 4500 23190 4860 23224
rect 5400 23276 5760 23310
rect 5400 23224 5429 23276
rect 5481 23224 5554 23276
rect 5606 23224 5679 23276
rect 5731 23224 5760 23276
rect 5400 23190 5760 23224
rect 6310 23276 6670 23310
rect 6310 23224 6339 23276
rect 6391 23224 6464 23276
rect 6516 23224 6589 23276
rect 6641 23224 6670 23276
rect 6310 23190 6670 23224
rect 6940 23276 7300 23310
rect 6940 23224 6969 23276
rect 7021 23224 7094 23276
rect 7146 23224 7219 23276
rect 7271 23224 7300 23276
rect 6940 23190 7300 23224
rect 8130 23276 8490 23310
rect 8130 23224 8159 23276
rect 8211 23224 8284 23276
rect 8336 23224 8409 23276
rect 8461 23224 8490 23276
rect 8130 23190 8490 23224
rect 9730 23276 10090 23310
rect 9730 23224 9759 23276
rect 9811 23224 9884 23276
rect 9936 23224 10009 23276
rect 10061 23224 10090 23276
rect 9730 23190 10090 23224
rect 11300 23276 11660 23310
rect 11300 23224 11329 23276
rect 11381 23224 11454 23276
rect 11506 23224 11579 23276
rect 11631 23224 11660 23276
rect 11300 23190 11660 23224
rect 13020 23276 13380 23310
rect 13020 23224 13049 23276
rect 13101 23224 13174 23276
rect 13226 23224 13299 23276
rect 13351 23224 13380 23276
rect 13020 23190 13380 23224
rect 15830 23266 16190 23300
rect 15830 23214 15859 23266
rect 15911 23214 15984 23266
rect 16036 23214 16109 23266
rect 16161 23214 16190 23266
rect -840 23100 -390 23129
rect 950 22680 1250 23180
rect 1830 22680 2130 23190
rect 2740 22680 3040 23190
rect 3620 22680 3920 23190
rect 4530 22680 4830 23190
rect 5430 22680 5730 23190
rect 6330 22680 6630 23190
rect 6940 22680 7240 23190
rect 8130 22680 8430 23190
rect 9730 22680 10030 23190
rect 11300 22680 11600 23190
rect 13020 22800 13320 23190
rect 15830 23180 16190 23214
rect 19390 23266 19750 23300
rect 19390 23214 19419 23266
rect 19471 23214 19544 23266
rect 19596 23214 19669 23266
rect 19721 23214 19750 23266
rect 19390 23180 19750 23214
rect 22670 23266 23030 23300
rect 22670 23214 22699 23266
rect 22751 23214 22824 23266
rect 22876 23214 22949 23266
rect 23001 23214 23030 23266
rect 22670 23180 23030 23214
rect 15830 22810 16130 23180
rect 19400 22810 19700 23180
rect 22670 22810 22920 23180
rect 12430 21360 13230 21670
rect 23210 19521 23330 19550
rect 23210 19480 23244 19521
rect 12500 19331 13240 19480
rect 12500 19279 12614 19331
rect 12666 19279 13240 19331
rect 12500 19206 13240 19279
rect 22900 19469 23244 19480
rect 23296 19490 23330 19521
rect 23296 19469 23340 19490
rect 22900 19396 23340 19469
rect 22900 19344 23244 19396
rect 23296 19344 23340 19396
rect 22900 19271 23340 19344
rect 12500 19154 12614 19206
rect 12666 19190 13240 19206
rect 12666 19154 12790 19190
rect 17110 19170 17970 19220
rect 22900 19219 23244 19271
rect 23296 19219 23340 19271
rect 22900 19190 23340 19219
rect 12500 19081 12790 19154
rect 12500 19029 12614 19081
rect 12666 19029 12790 19081
rect 12500 18750 12790 19029
rect 17430 18830 17510 19170
rect 17880 18870 17970 19170
rect 17110 18750 17510 18830
rect 12500 18670 12810 18750
rect 17430 18670 17510 18750
rect 12500 18660 12820 18670
rect 12500 18601 12890 18660
rect 12500 18549 12614 18601
rect 12666 18549 12890 18601
rect 13130 18590 13340 18670
rect 10780 18356 11330 18490
rect 10780 18304 11079 18356
rect 11131 18304 11204 18356
rect 11256 18304 11330 18356
rect 10780 18190 11330 18304
rect 12500 18476 12890 18549
rect 12500 18424 12614 18476
rect 12666 18424 12890 18476
rect 12500 18351 12890 18424
rect 12500 18299 12614 18351
rect 12666 18299 12890 18351
rect 12500 18130 12890 18299
rect 13140 18130 13240 18590
rect 17110 18330 17510 18670
rect 17890 18330 17970 18870
rect 23070 18750 23300 19190
rect 23450 19036 23550 19060
rect 23450 18984 23474 19036
rect 23526 18984 23550 19036
rect 15020 16456 15180 16470
rect 15020 16404 15034 16456
rect 15086 16404 15114 16456
rect 15166 16404 15180 16456
rect 15020 16390 15180 16404
rect 14500 16346 14680 16360
rect 14500 16294 14514 16346
rect 14566 16294 14614 16346
rect 14666 16294 14680 16346
rect 14500 16280 14680 16294
rect 14580 16166 14680 16280
rect 14580 16114 14604 16166
rect 14656 16114 14680 16166
rect 14580 16046 14680 16114
rect 14580 15994 14604 16046
rect 14656 15994 14680 16046
rect 870 14986 1230 15020
rect 870 14934 899 14986
rect 951 14934 1024 14986
rect 1076 14934 1149 14986
rect 1201 14934 1230 14986
rect 870 14866 1230 14934
rect 870 14814 899 14866
rect 951 14814 1024 14866
rect 1076 14814 1149 14866
rect 1201 14814 1230 14866
rect 870 13670 1230 14814
rect 2590 14986 2950 15020
rect 2590 14934 2619 14986
rect 2671 14934 2744 14986
rect 2796 14934 2869 14986
rect 2921 14934 2950 14986
rect 2590 14866 2950 14934
rect 2590 14814 2619 14866
rect 2671 14814 2744 14866
rect 2796 14814 2869 14866
rect 2921 14814 2950 14866
rect 2590 13670 2950 14814
rect 4030 14986 4390 15020
rect 4030 14934 4059 14986
rect 4111 14934 4184 14986
rect 4236 14934 4309 14986
rect 4361 14934 4390 14986
rect 4030 14866 4390 14934
rect 4030 14814 4059 14866
rect 4111 14814 4184 14866
rect 4236 14814 4309 14866
rect 4361 14814 4390 14866
rect 4030 13670 4390 14814
rect 5490 14986 5850 15020
rect 5490 14934 5519 14986
rect 5571 14934 5644 14986
rect 5696 14934 5769 14986
rect 5821 14934 5850 14986
rect 5490 14866 5850 14934
rect 5490 14814 5519 14866
rect 5571 14814 5644 14866
rect 5696 14814 5769 14866
rect 5821 14814 5850 14866
rect 5490 13670 5850 14814
rect 7330 14946 7690 14980
rect 7330 14894 7359 14946
rect 7411 14894 7484 14946
rect 7536 14894 7609 14946
rect 7661 14894 7690 14946
rect 7330 13670 7690 14894
rect 8800 14956 9160 14990
rect 8800 14904 8829 14956
rect 8881 14904 8954 14956
rect 9006 14904 9079 14956
rect 9131 14904 9160 14956
rect -7000 12906 -6900 12930
rect -7000 12854 -6976 12906
rect -6924 12854 -6900 12906
rect -7000 12830 -6900 12854
rect -7370 12766 -7270 12790
rect -7370 12714 -7346 12766
rect -7294 12714 -7270 12766
rect -7370 12690 -7270 12714
rect -7650 12686 -7570 12690
rect -7650 12634 -7636 12686
rect -7584 12634 -7570 12686
rect -7650 12630 -7570 12634
rect -8550 12596 -8470 12600
rect -8550 12544 -8536 12596
rect -8484 12544 -8470 12596
rect -8550 12540 -8470 12544
rect -9450 12476 -9370 12480
rect -9450 12424 -9436 12476
rect -9384 12424 -9370 12476
rect -9450 12420 -9370 12424
rect -9750 12296 -9670 12300
rect -9750 12244 -9736 12296
rect -9684 12244 -9670 12296
rect -9450 12270 -9390 12420
rect -9150 12386 -9070 12390
rect -9150 12334 -9136 12386
rect -9084 12334 -9070 12386
rect -9150 12330 -9070 12334
rect -9130 12270 -9070 12330
rect -8850 12386 -8770 12390
rect -8850 12334 -8836 12386
rect -8784 12334 -8770 12386
rect -8850 12330 -8770 12334
rect -9750 12240 -9670 12244
rect -8850 12240 -8790 12330
rect -8530 12260 -8470 12540
rect -8250 12296 -8170 12300
rect -8250 12244 -8236 12296
rect -8184 12244 -8170 12296
rect -8250 12240 -8170 12244
rect -7630 12240 -7570 12630
rect -7330 12240 -7270 12690
rect -7940 12206 -7870 12210
rect -7940 12154 -7936 12206
rect -7884 12154 -7870 12206
rect -7940 12150 -7870 12154
rect -6980 11680 -6900 12830
rect -6480 11480 -6380 13140
rect 8800 12840 9160 14904
rect 11660 14966 12020 15000
rect 11660 14914 11689 14966
rect 11741 14914 11814 14966
rect 11866 14914 11939 14966
rect 11991 14914 12020 14966
rect 11660 14880 12020 14914
rect 12670 14966 13030 15000
rect 12670 14914 12699 14966
rect 12751 14914 12824 14966
rect 12876 14914 12949 14966
rect 13001 14914 13030 14966
rect 12670 14880 13030 14914
rect 14580 14956 14680 15994
rect 14580 14904 14604 14956
rect 14656 14904 14680 14956
rect 14580 14890 14680 14904
rect 15080 15906 15180 16390
rect 15080 15854 15104 15906
rect 15156 15854 15180 15906
rect 15080 15786 15180 15854
rect 15080 15734 15104 15786
rect 15156 15734 15180 15786
rect 11680 14700 12000 14880
rect 12700 14730 13000 14880
rect 15080 14846 15180 15734
rect 20270 16346 20350 16360
rect 20270 16294 20284 16346
rect 20336 16294 20350 16346
rect 15080 14794 15104 14846
rect 15156 14794 15180 14846
rect 15080 14780 15180 14794
rect 15240 14966 15600 15000
rect 15240 14914 15269 14966
rect 15321 14914 15394 14966
rect 15446 14914 15519 14966
rect 15571 14914 15600 14966
rect 15240 14880 15600 14914
rect 15720 14966 16080 15000
rect 15720 14914 15749 14966
rect 15801 14914 15874 14966
rect 15926 14914 15999 14966
rect 16051 14914 16080 14966
rect 15720 14880 16080 14914
rect 15240 14730 15500 14880
rect 15720 14430 15940 14880
rect 20270 14550 20350 16294
rect 20390 16346 20470 16360
rect 20390 16294 20404 16346
rect 20456 16294 20470 16346
rect 20390 14646 20470 16294
rect 22280 16336 22400 16350
rect 22280 16284 22314 16336
rect 22366 16284 22400 16336
rect 20390 14594 20404 14646
rect 20456 14594 20470 14646
rect 20390 14580 20470 14594
rect 20500 14946 21220 14980
rect 20500 14894 20529 14946
rect 20581 14894 20654 14946
rect 20706 14894 20779 14946
rect 20831 14894 20889 14946
rect 20941 14894 21014 14946
rect 21066 14894 21139 14946
rect 21191 14894 21220 14946
rect 20500 14860 21220 14894
rect 20250 14526 20350 14550
rect 20250 14474 20274 14526
rect 20326 14474 20350 14526
rect 20250 14460 20350 14474
rect 20500 14430 20700 14860
rect 15940 14320 16100 14420
rect 20410 14230 20700 14430
rect 20810 14430 21220 14860
rect 20810 14320 21260 14430
rect 22280 14196 22400 16284
rect 23450 14406 23550 18984
rect 23690 16496 23890 16520
rect 23690 16444 23714 16496
rect 23766 16444 23814 16496
rect 23866 16444 23890 16496
rect 23690 16420 23890 16444
rect 29662 16270 29742 16320
rect 29500 16190 29742 16270
rect 29500 16166 29600 16190
rect 29500 16114 29524 16166
rect 29576 16114 29600 16166
rect 29500 16086 29600 16114
rect 29500 16034 29524 16086
rect 29576 16034 29600 16086
rect 29500 16010 29600 16034
rect 29320 15906 29420 15930
rect 29320 15854 29344 15906
rect 29396 15854 29420 15906
rect 29320 15826 29420 15854
rect 29320 15774 29344 15826
rect 29396 15774 29420 15826
rect 29320 15750 29420 15774
rect 23450 14354 23474 14406
rect 23526 14354 23550 14406
rect 23450 14340 23550 14354
rect 22280 14144 22314 14196
rect 22366 14144 22400 14196
rect 22280 14120 22400 14144
rect 20780 12930 21200 12940
rect 16310 12750 16610 12760
rect -6710 11456 -6380 11480
rect -6710 11404 -6576 11456
rect -6524 11404 -6456 11456
rect -6404 11404 -6380 11456
rect -6710 11380 -6380 11404
rect 14120 10870 14430 12650
rect 15240 11680 15550 12710
rect 16310 11670 16620 12750
rect 19660 11660 19960 12750
rect 20260 12730 21200 12930
rect 20500 12700 21200 12730
rect 20500 11520 20800 12700
rect 21340 11660 21640 12710
rect 900 7476 1200 7610
rect 900 7424 959 7476
rect 1011 7424 1084 7476
rect 1136 7424 1200 7476
rect 900 7300 1200 7424
rect 1510 7476 1810 7630
rect 1510 7424 1569 7476
rect 1621 7424 1694 7476
rect 1746 7424 1810 7476
rect 1510 7280 1810 7424
rect 2660 7476 2960 7630
rect 2660 7424 2719 7476
rect 2771 7424 2844 7476
rect 2896 7424 2960 7476
rect 2660 7280 2960 7424
rect 3830 7476 4130 7630
rect 3830 7424 3889 7476
rect 3941 7424 4014 7476
rect 4066 7424 4130 7476
rect 3830 7280 4130 7424
rect 4990 7476 5290 7630
rect 4990 7424 5049 7476
rect 5101 7424 5174 7476
rect 5226 7424 5290 7476
rect 4990 7280 5290 7424
rect 6160 7476 6450 7630
rect 6160 7424 6219 7476
rect 6271 7424 6344 7476
rect 6396 7424 6450 7476
rect 6160 7280 6450 7424
rect 7320 7476 7620 7630
rect 7320 7424 7379 7476
rect 7431 7424 7504 7476
rect 7556 7424 7620 7476
rect 7320 7300 7620 7424
rect 1370 406 1730 560
rect 1370 354 1399 406
rect 1451 354 1524 406
rect 1576 354 1649 406
rect 1701 354 1730 406
rect 1370 320 1730 354
rect 3100 406 3460 560
rect 3100 354 3129 406
rect 3181 354 3254 406
rect 3306 354 3379 406
rect 3431 354 3460 406
rect 3100 320 3460 354
rect 5160 406 5520 560
rect 5160 354 5189 406
rect 5241 354 5314 406
rect 5366 354 5439 406
rect 5491 354 5520 406
rect 5160 320 5520 354
rect 8800 396 9160 560
rect 8800 344 8829 396
rect 8881 344 8954 396
rect 9006 344 9079 396
rect 9131 344 9160 396
rect 8800 310 9160 344
rect 10920 396 11280 560
rect 10920 344 10949 396
rect 11001 344 11074 396
rect 11126 344 11199 396
rect 11251 344 11280 396
rect 10920 310 11280 344
rect 14650 396 15010 560
rect 14650 344 14679 396
rect 14731 344 14804 396
rect 14856 344 14929 396
rect 14981 344 15010 396
rect 14650 310 15010 344
rect 17010 396 17370 560
rect 17010 344 17039 396
rect 17091 344 17164 396
rect 17216 344 17289 396
rect 17341 344 17370 396
rect 17010 310 17370 344
rect 19020 396 19380 560
rect 19020 344 19049 396
rect 19101 344 19174 396
rect 19226 344 19299 396
rect 19351 344 19380 396
rect 19020 310 19380 344
rect 20980 396 21340 430
rect 20980 344 21009 396
rect 21061 344 21134 396
rect 21186 344 21259 396
rect 21311 344 21340 396
rect 20980 310 21340 344
<< via1 >>
rect -10411 25214 -10359 25266
rect -10286 25214 -10234 25266
rect -10161 25214 -10109 25266
rect -8641 25224 -8589 25276
rect -8516 25224 -8464 25276
rect -8391 25224 -8339 25276
rect -6911 25214 -6859 25266
rect -6786 25214 -6734 25266
rect -6661 25214 -6609 25266
rect -466 24569 -414 24621
rect -466 24444 -414 24496
rect -466 24319 -414 24371
rect -486 23379 -434 23431
rect -486 23254 -434 23306
rect -486 23129 -434 23181
rect 969 23214 1021 23266
rect 1094 23214 1146 23266
rect 1219 23214 1271 23266
rect 1839 23224 1891 23276
rect 1964 23224 2016 23276
rect 2089 23224 2141 23276
rect 2739 23224 2791 23276
rect 2864 23224 2916 23276
rect 2989 23224 3041 23276
rect 3639 23224 3691 23276
rect 3764 23224 3816 23276
rect 3889 23224 3941 23276
rect 4529 23224 4581 23276
rect 4654 23224 4706 23276
rect 4779 23224 4831 23276
rect 5429 23224 5481 23276
rect 5554 23224 5606 23276
rect 5679 23224 5731 23276
rect 6339 23224 6391 23276
rect 6464 23224 6516 23276
rect 6589 23224 6641 23276
rect 6969 23224 7021 23276
rect 7094 23224 7146 23276
rect 7219 23224 7271 23276
rect 8159 23224 8211 23276
rect 8284 23224 8336 23276
rect 8409 23224 8461 23276
rect 9759 23224 9811 23276
rect 9884 23224 9936 23276
rect 10009 23224 10061 23276
rect 11329 23224 11381 23276
rect 11454 23224 11506 23276
rect 11579 23224 11631 23276
rect 13049 23224 13101 23276
rect 13174 23224 13226 23276
rect 13299 23224 13351 23276
rect 15859 23214 15911 23266
rect 15984 23214 16036 23266
rect 16109 23214 16161 23266
rect 19419 23214 19471 23266
rect 19544 23214 19596 23266
rect 19669 23214 19721 23266
rect 22699 23214 22751 23266
rect 22824 23214 22876 23266
rect 22949 23214 23001 23266
rect 12614 19279 12666 19331
rect 23244 19469 23296 19521
rect 23244 19344 23296 19396
rect 12614 19154 12666 19206
rect 23244 19219 23296 19271
rect 12614 19029 12666 19081
rect 12614 18549 12666 18601
rect 11079 18304 11131 18356
rect 11204 18304 11256 18356
rect 12614 18424 12666 18476
rect 12614 18299 12666 18351
rect 23474 18984 23526 19036
rect 15034 16404 15086 16456
rect 15114 16404 15166 16456
rect 14514 16294 14566 16346
rect 14614 16294 14666 16346
rect 14604 16114 14656 16166
rect 14604 15994 14656 16046
rect 899 14934 951 14986
rect 1024 14934 1076 14986
rect 1149 14934 1201 14986
rect 899 14814 951 14866
rect 1024 14814 1076 14866
rect 1149 14814 1201 14866
rect 2619 14934 2671 14986
rect 2744 14934 2796 14986
rect 2869 14934 2921 14986
rect 2619 14814 2671 14866
rect 2744 14814 2796 14866
rect 2869 14814 2921 14866
rect 4059 14934 4111 14986
rect 4184 14934 4236 14986
rect 4309 14934 4361 14986
rect 4059 14814 4111 14866
rect 4184 14814 4236 14866
rect 4309 14814 4361 14866
rect 5519 14934 5571 14986
rect 5644 14934 5696 14986
rect 5769 14934 5821 14986
rect 5519 14814 5571 14866
rect 5644 14814 5696 14866
rect 5769 14814 5821 14866
rect 7359 14894 7411 14946
rect 7484 14894 7536 14946
rect 7609 14894 7661 14946
rect 8829 14904 8881 14956
rect 8954 14904 9006 14956
rect 9079 14904 9131 14956
rect -6976 12854 -6924 12906
rect -7346 12714 -7294 12766
rect -7636 12634 -7584 12686
rect -8536 12544 -8484 12596
rect -9436 12424 -9384 12476
rect -9736 12244 -9684 12296
rect -9136 12334 -9084 12386
rect -8836 12334 -8784 12386
rect -8236 12244 -8184 12296
rect -7936 12154 -7884 12206
rect 11689 14914 11741 14966
rect 11814 14914 11866 14966
rect 11939 14914 11991 14966
rect 12699 14914 12751 14966
rect 12824 14914 12876 14966
rect 12949 14914 13001 14966
rect 14604 14904 14656 14956
rect 15104 15854 15156 15906
rect 15104 15734 15156 15786
rect 20284 16294 20336 16346
rect 15104 14794 15156 14846
rect 15269 14914 15321 14966
rect 15394 14914 15446 14966
rect 15519 14914 15571 14966
rect 15749 14914 15801 14966
rect 15874 14914 15926 14966
rect 15999 14914 16051 14966
rect 20404 16294 20456 16346
rect 22314 16284 22366 16336
rect 20404 14594 20456 14646
rect 20529 14894 20581 14946
rect 20654 14894 20706 14946
rect 20779 14894 20831 14946
rect 20889 14894 20941 14946
rect 21014 14894 21066 14946
rect 21139 14894 21191 14946
rect 20274 14474 20326 14526
rect 23714 16444 23766 16496
rect 23814 16444 23866 16496
rect 29524 16114 29576 16166
rect 29524 16034 29576 16086
rect 29344 15854 29396 15906
rect 29344 15774 29396 15826
rect 23474 14354 23526 14406
rect 22314 14144 22366 14196
rect -6576 11404 -6524 11456
rect -6456 11404 -6404 11456
rect 959 7424 1011 7476
rect 1084 7424 1136 7476
rect 1569 7424 1621 7476
rect 1694 7424 1746 7476
rect 2719 7424 2771 7476
rect 2844 7424 2896 7476
rect 3889 7424 3941 7476
rect 4014 7424 4066 7476
rect 5049 7424 5101 7476
rect 5174 7424 5226 7476
rect 6219 7424 6271 7476
rect 6344 7424 6396 7476
rect 7379 7424 7431 7476
rect 7504 7424 7556 7476
rect 1399 354 1451 406
rect 1524 354 1576 406
rect 1649 354 1701 406
rect 3129 354 3181 406
rect 3254 354 3306 406
rect 3379 354 3431 406
rect 5189 354 5241 406
rect 5314 354 5366 406
rect 5439 354 5491 406
rect 8829 344 8881 396
rect 8954 344 9006 396
rect 9079 344 9131 396
rect 10949 344 11001 396
rect 11074 344 11126 396
rect 11199 344 11251 396
rect 14679 344 14731 396
rect 14804 344 14856 396
rect 14929 344 14981 396
rect 17039 344 17091 396
rect 17164 344 17216 396
rect 17289 344 17341 396
rect 19049 344 19101 396
rect 19174 344 19226 396
rect 19299 344 19351 396
rect 21009 344 21061 396
rect 21134 344 21186 396
rect 21259 344 21311 396
<< metal2 >>
rect -10440 25268 -10080 25300
rect -10440 25212 -10413 25268
rect -10357 25212 -10288 25268
rect -10232 25212 -10163 25268
rect -10107 25212 -10080 25268
rect -10440 25180 -10080 25212
rect -8670 25278 -8310 25310
rect -8670 25222 -8643 25278
rect -8587 25222 -8518 25278
rect -8462 25222 -8393 25278
rect -8337 25222 -8310 25278
rect -8670 25190 -8310 25222
rect -6940 25268 -6580 25300
rect -6940 25212 -6913 25268
rect -6857 25212 -6788 25268
rect -6732 25212 -6663 25268
rect -6607 25212 -6580 25268
rect -6940 25180 -6580 25212
rect -500 24623 -380 24650
rect -500 24567 -468 24623
rect -412 24567 -380 24623
rect -500 24498 -380 24567
rect -500 24442 -468 24498
rect -412 24442 -380 24498
rect -500 24373 -380 24442
rect -500 24317 -468 24373
rect -412 24317 -380 24373
rect -500 24290 -380 24317
rect -520 23433 -400 23460
rect -520 23377 -488 23433
rect -432 23377 -400 23433
rect -520 23308 -400 23377
rect -520 23252 -488 23308
rect -432 23252 -400 23308
rect -520 23183 -400 23252
rect -520 23127 -488 23183
rect -432 23127 -400 23183
rect 940 23268 1300 23300
rect 940 23212 967 23268
rect 1023 23212 1092 23268
rect 1148 23212 1217 23268
rect 1273 23212 1300 23268
rect 940 23180 1300 23212
rect 1810 23278 2170 23310
rect 1810 23222 1837 23278
rect 1893 23222 1962 23278
rect 2018 23222 2087 23278
rect 2143 23222 2170 23278
rect 1810 23190 2170 23222
rect 2710 23278 3070 23310
rect 2710 23222 2737 23278
rect 2793 23222 2862 23278
rect 2918 23222 2987 23278
rect 3043 23222 3070 23278
rect 2710 23190 3070 23222
rect 3610 23278 3970 23310
rect 3610 23222 3637 23278
rect 3693 23222 3762 23278
rect 3818 23222 3887 23278
rect 3943 23222 3970 23278
rect 3610 23190 3970 23222
rect 4500 23278 4860 23310
rect 4500 23222 4527 23278
rect 4583 23222 4652 23278
rect 4708 23222 4777 23278
rect 4833 23222 4860 23278
rect 4500 23190 4860 23222
rect 5400 23278 5760 23310
rect 5400 23222 5427 23278
rect 5483 23222 5552 23278
rect 5608 23222 5677 23278
rect 5733 23222 5760 23278
rect 5400 23190 5760 23222
rect 6310 23278 6670 23310
rect 6310 23222 6337 23278
rect 6393 23222 6462 23278
rect 6518 23222 6587 23278
rect 6643 23222 6670 23278
rect 6310 23190 6670 23222
rect 6940 23278 7300 23310
rect 6940 23222 6967 23278
rect 7023 23222 7092 23278
rect 7148 23222 7217 23278
rect 7273 23222 7300 23278
rect 6940 23190 7300 23222
rect 8130 23278 8490 23310
rect 8130 23222 8157 23278
rect 8213 23222 8282 23278
rect 8338 23222 8407 23278
rect 8463 23222 8490 23278
rect 8130 23190 8490 23222
rect 9730 23278 10090 23310
rect 9730 23222 9757 23278
rect 9813 23222 9882 23278
rect 9938 23222 10007 23278
rect 10063 23222 10090 23278
rect 9730 23190 10090 23222
rect 11300 23278 11660 23310
rect 11300 23222 11327 23278
rect 11383 23222 11452 23278
rect 11508 23222 11577 23278
rect 11633 23222 11660 23278
rect 11300 23190 11660 23222
rect 13020 23278 13380 23310
rect 13020 23222 13047 23278
rect 13103 23222 13172 23278
rect 13228 23222 13297 23278
rect 13353 23222 13380 23278
rect 13020 23190 13380 23222
rect 15830 23268 16190 23300
rect 15830 23212 15857 23268
rect 15913 23212 15982 23268
rect 16038 23212 16107 23268
rect 16163 23212 16190 23268
rect 15830 23180 16190 23212
rect 19390 23268 19750 23300
rect 19390 23212 19417 23268
rect 19473 23212 19542 23268
rect 19598 23212 19667 23268
rect 19723 23212 19750 23268
rect 19390 23180 19750 23212
rect 22670 23268 23030 23300
rect 22670 23212 22697 23268
rect 22753 23212 22822 23268
rect 22878 23212 22947 23268
rect 23003 23212 23030 23268
rect 22670 23180 23030 23212
rect -520 23100 -400 23127
rect 23210 19523 23330 19550
rect 23210 19467 23242 19523
rect 23298 19467 23330 19523
rect 23210 19398 23330 19467
rect 12580 19333 12700 19360
rect 12580 19277 12612 19333
rect 12668 19277 12700 19333
rect 12580 19208 12700 19277
rect 12580 19152 12612 19208
rect 12668 19152 12700 19208
rect 23210 19342 23242 19398
rect 23298 19342 23330 19398
rect 23210 19273 23330 19342
rect 23210 19217 23242 19273
rect 23298 19217 23330 19273
rect 23210 19190 23330 19217
rect 12580 19083 12700 19152
rect 12580 19027 12612 19083
rect 12668 19027 12700 19083
rect 12580 19000 12700 19027
rect 23070 19038 23550 19060
rect 23070 18982 23087 19038
rect 23143 19036 23550 19038
rect 23143 18984 23474 19036
rect 23526 18984 23550 19036
rect 23143 18982 23550 18984
rect 23070 18960 23550 18982
rect 12580 18603 12700 18630
rect 12580 18547 12612 18603
rect 12668 18547 12700 18603
rect 12580 18478 12700 18547
rect 12580 18422 12612 18478
rect 12668 18422 12700 18478
rect 11050 18358 11290 18390
rect 11050 18302 11077 18358
rect 11133 18302 11202 18358
rect 11258 18302 11290 18358
rect 11050 18270 11290 18302
rect 12580 18353 12700 18422
rect 12580 18297 12612 18353
rect 12668 18297 12700 18353
rect 12580 18270 12700 18297
rect 23690 16498 23890 16520
rect 15020 16460 15110 16470
rect 15020 16456 15170 16460
rect 15020 16404 15034 16456
rect 15086 16404 15114 16456
rect 15166 16404 15170 16456
rect 23690 16442 23712 16498
rect 23768 16442 23812 16498
rect 23868 16442 23890 16498
rect 23690 16420 23890 16442
rect 15020 16400 15170 16404
rect 15020 16390 15110 16400
rect 14500 16348 14580 16360
rect 14500 16292 14512 16348
rect 14568 16292 14580 16348
rect 14500 16280 14580 16292
rect 14590 16348 14670 16350
rect 14590 16292 14612 16348
rect 14668 16292 14670 16348
rect 14590 16290 14670 16292
rect 20280 16346 20340 16350
rect 20280 16294 20284 16346
rect 20336 16294 20340 16346
rect 20280 16290 20340 16294
rect 20390 16346 20470 16360
rect 20390 16294 20404 16346
rect 20456 16294 20470 16346
rect 20390 16280 20470 16294
rect 22280 16338 22400 16350
rect 22280 16282 22312 16338
rect 22368 16282 22400 16338
rect 22280 16270 22400 16282
rect 29320 16320 29590 16410
rect 14580 16168 14680 16190
rect 14580 16112 14602 16168
rect 14658 16112 14680 16168
rect 14580 16048 14680 16112
rect 14580 15992 14602 16048
rect 14658 15992 14680 16048
rect 14580 15970 14680 15992
rect 15080 15908 15180 15930
rect 15080 15852 15102 15908
rect 15158 15852 15180 15908
rect 15080 15788 15180 15852
rect 15080 15732 15102 15788
rect 15158 15732 15180 15788
rect 29320 15908 29420 16320
rect 29500 16168 29600 16190
rect 29500 16112 29522 16168
rect 29578 16112 29600 16168
rect 29500 16088 29600 16112
rect 29500 16032 29522 16088
rect 29578 16032 29600 16088
rect 29500 16010 29600 16032
rect 29320 15852 29342 15908
rect 29398 15852 29420 15908
rect 29320 15828 29420 15852
rect 29320 15772 29342 15828
rect 29398 15772 29420 15828
rect 29320 15750 29420 15772
rect 15080 15710 15180 15732
rect 870 14988 1230 15020
rect 870 14932 897 14988
rect 953 14932 1022 14988
rect 1078 14932 1147 14988
rect 1203 14932 1230 14988
rect 870 14868 1230 14932
rect 870 14812 897 14868
rect 953 14812 1022 14868
rect 1078 14812 1147 14868
rect 1203 14812 1230 14868
rect 870 14780 1230 14812
rect 2590 14988 2950 15020
rect 2590 14932 2617 14988
rect 2673 14932 2742 14988
rect 2798 14932 2867 14988
rect 2923 14932 2950 14988
rect 2590 14868 2950 14932
rect 2590 14812 2617 14868
rect 2673 14812 2742 14868
rect 2798 14812 2867 14868
rect 2923 14812 2950 14868
rect 2590 14780 2950 14812
rect 4030 14988 4390 15020
rect 4030 14932 4057 14988
rect 4113 14932 4182 14988
rect 4238 14932 4307 14988
rect 4363 14932 4390 14988
rect 4030 14868 4390 14932
rect 4030 14812 4057 14868
rect 4113 14812 4182 14868
rect 4238 14812 4307 14868
rect 4363 14812 4390 14868
rect 4030 14780 4390 14812
rect 5490 14988 5850 15020
rect 5490 14932 5517 14988
rect 5573 14932 5642 14988
rect 5698 14932 5767 14988
rect 5823 14932 5850 14988
rect 5490 14868 5850 14932
rect 5490 14812 5517 14868
rect 5573 14812 5642 14868
rect 5698 14812 5767 14868
rect 5823 14812 5850 14868
rect 7330 14948 7690 14980
rect 7330 14892 7357 14948
rect 7413 14892 7482 14948
rect 7538 14892 7607 14948
rect 7663 14892 7690 14948
rect 7330 14860 7690 14892
rect 8800 14958 9160 14990
rect 8800 14902 8827 14958
rect 8883 14902 8952 14958
rect 9008 14902 9077 14958
rect 9133 14902 9160 14958
rect 8800 14870 9160 14902
rect 11660 14968 12020 15000
rect 11660 14912 11687 14968
rect 11743 14912 11812 14968
rect 11868 14912 11937 14968
rect 11993 14912 12020 14968
rect 11660 14880 12020 14912
rect 12670 14968 13030 15000
rect 12670 14912 12697 14968
rect 12753 14912 12822 14968
rect 12878 14912 12947 14968
rect 13003 14912 13030 14968
rect 12670 14880 13030 14912
rect 14580 14958 14680 14970
rect 14580 14902 14602 14958
rect 14658 14902 14680 14958
rect 14580 14890 14680 14902
rect 15240 14968 15600 15000
rect 15240 14912 15267 14968
rect 15323 14912 15392 14968
rect 15448 14912 15517 14968
rect 15573 14912 15600 14968
rect 15240 14880 15600 14912
rect 15720 14968 16080 15000
rect 15720 14912 15747 14968
rect 15803 14912 15872 14968
rect 15928 14912 15997 14968
rect 16053 14912 16080 14968
rect 15720 14880 16080 14912
rect 20500 14948 21220 14980
rect 20500 14892 20527 14948
rect 20583 14892 20652 14948
rect 20708 14892 20777 14948
rect 20833 14892 20887 14948
rect 20943 14892 21012 14948
rect 21068 14892 21137 14948
rect 21193 14892 21220 14948
rect 20500 14860 21220 14892
rect 5490 14780 5850 14812
rect 15090 14846 15170 14850
rect 15090 14794 15104 14846
rect 15156 14794 15170 14846
rect 15090 14790 15170 14794
rect 15960 14646 20470 14660
rect 15960 14594 20404 14646
rect 20456 14594 20470 14646
rect 15960 14580 20470 14594
rect 16070 14528 16170 14550
rect 16070 14472 16092 14528
rect 16148 14472 16170 14528
rect 16070 14450 16170 14472
rect 20250 14528 20350 14550
rect 20250 14472 20272 14528
rect 20328 14472 20350 14528
rect 20250 14460 20350 14472
rect 21130 14406 23550 14420
rect 21130 14354 23474 14406
rect 23526 14354 23550 14406
rect 21130 14340 23550 14354
rect 21130 14290 21210 14340
rect 22280 14198 22400 14220
rect 22280 14142 22312 14198
rect 22368 14142 22400 14198
rect 22280 14120 22400 14142
rect 21240 14058 21320 14070
rect 21240 14002 21252 14058
rect 21308 14002 21320 14058
rect 21240 13990 21320 14002
rect -7000 12908 -6900 12930
rect -7000 12852 -6978 12908
rect -6922 12852 -6900 12908
rect -7000 12830 -6900 12852
rect -7370 12768 -7270 12790
rect -7370 12712 -7348 12768
rect -7292 12712 -7270 12768
rect -10890 12698 -10810 12710
rect -10890 12642 -10878 12698
rect -10822 12690 -10810 12698
rect -7370 12690 -7270 12712
rect -10822 12686 -7570 12690
rect -10822 12642 -7636 12686
rect -10890 12634 -7636 12642
rect -7584 12634 -7570 12686
rect -10890 12630 -7570 12634
rect -10750 12596 -8470 12600
rect -10750 12588 -8536 12596
rect -10750 12532 -10738 12588
rect -10682 12544 -8536 12588
rect -8484 12544 -8470 12596
rect -10682 12540 -8470 12544
rect -10682 12532 -10670 12540
rect -10750 12520 -10670 12532
rect -5930 12480 -5850 13200
rect -9450 12476 -5850 12480
rect -9450 12424 -9436 12476
rect -9384 12424 -5850 12476
rect -9450 12420 -5850 12424
rect -10470 12398 -10390 12410
rect -10470 12342 -10458 12398
rect -10402 12390 -10390 12398
rect -5820 12390 -5740 13010
rect -10402 12386 -9070 12390
rect -10402 12342 -9136 12386
rect -10470 12334 -9136 12342
rect -9084 12334 -9070 12386
rect -10470 12330 -9070 12334
rect -8850 12386 -5740 12390
rect -8850 12334 -8836 12386
rect -8784 12334 -5740 12386
rect -8850 12330 -5740 12334
rect -5710 12300 -5630 13010
rect -10330 12296 -9670 12300
rect -10330 12288 -9736 12296
rect -10330 12232 -10318 12288
rect -10262 12244 -9736 12288
rect -9684 12244 -9670 12296
rect -10262 12240 -9670 12244
rect -8250 12296 -5630 12300
rect -8250 12244 -8236 12296
rect -8184 12244 -5630 12296
rect -8250 12240 -5630 12244
rect -10262 12232 -10250 12240
rect -10330 12220 -10250 12232
rect -5600 12210 -5520 13370
rect -7950 12206 -5520 12210
rect -7950 12154 -7936 12206
rect -7884 12154 -5520 12206
rect -7950 12150 -5520 12154
rect -10090 12060 -9860 12120
rect -6630 12103 -5990 12120
rect -6630 12060 -6148 12103
rect -6170 12047 -6148 12060
rect -6092 12047 -6058 12103
rect -6002 12047 -5990 12103
rect -6170 12020 -5990 12047
rect -10090 11940 -9870 12000
rect -6620 11880 -6560 12000
rect -6620 11863 -6190 11880
rect -6620 11820 -6358 11863
rect -6380 11807 -6358 11820
rect -6302 11807 -6268 11863
rect -6212 11820 -6190 11863
rect -6212 11807 -6200 11820
rect -6380 11780 -6200 11807
rect -6600 11458 -6380 11480
rect -6600 11402 -6578 11458
rect -6522 11402 -6458 11458
rect -6402 11402 -6380 11458
rect -6600 11380 -6380 11402
rect 930 7478 1170 7510
rect 930 7422 957 7478
rect 1013 7422 1082 7478
rect 1138 7422 1170 7478
rect 930 7390 1170 7422
rect 1540 7478 1780 7510
rect 1540 7422 1567 7478
rect 1623 7422 1692 7478
rect 1748 7422 1780 7478
rect 1540 7390 1780 7422
rect 2690 7478 2930 7510
rect 2690 7422 2717 7478
rect 2773 7422 2842 7478
rect 2898 7422 2930 7478
rect 2690 7390 2930 7422
rect 3860 7478 4100 7510
rect 3860 7422 3887 7478
rect 3943 7422 4012 7478
rect 4068 7422 4100 7478
rect 3860 7390 4100 7422
rect 5020 7478 5260 7510
rect 5020 7422 5047 7478
rect 5103 7422 5172 7478
rect 5228 7422 5260 7478
rect 5020 7390 5260 7422
rect 6190 7478 6430 7510
rect 6190 7422 6217 7478
rect 6273 7422 6342 7478
rect 6398 7422 6430 7478
rect 6190 7390 6430 7422
rect 7350 7478 7590 7510
rect 7350 7422 7377 7478
rect 7433 7422 7502 7478
rect 7558 7422 7590 7478
rect 7350 7390 7590 7422
rect 1370 408 1730 440
rect 1370 352 1397 408
rect 1453 352 1522 408
rect 1578 352 1647 408
rect 1703 352 1730 408
rect 1370 320 1730 352
rect 3100 408 3460 440
rect 3100 352 3127 408
rect 3183 352 3252 408
rect 3308 352 3377 408
rect 3433 352 3460 408
rect 3100 320 3460 352
rect 5160 408 5520 440
rect 5160 352 5187 408
rect 5243 352 5312 408
rect 5368 352 5437 408
rect 5493 352 5520 408
rect 5160 320 5520 352
rect 8800 398 9160 430
rect 8800 342 8827 398
rect 8883 342 8952 398
rect 9008 342 9077 398
rect 9133 342 9160 398
rect 8800 310 9160 342
rect 10920 398 11280 430
rect 10920 342 10947 398
rect 11003 342 11072 398
rect 11128 342 11197 398
rect 11253 342 11280 398
rect 10920 310 11280 342
rect 14650 398 15010 430
rect 14650 342 14677 398
rect 14733 342 14802 398
rect 14858 342 14927 398
rect 14983 342 15010 398
rect 14650 310 15010 342
rect 17010 398 17370 430
rect 17010 342 17037 398
rect 17093 342 17162 398
rect 17218 342 17287 398
rect 17343 342 17370 398
rect 17010 310 17370 342
rect 19020 398 19380 430
rect 19020 342 19047 398
rect 19103 342 19172 398
rect 19228 342 19297 398
rect 19353 342 19380 398
rect 19020 310 19380 342
rect 20980 398 21340 560
rect 20980 342 21007 398
rect 21063 342 21132 398
rect 21188 342 21257 398
rect 21313 342 21340 398
rect 20980 310 21340 342
<< via2 >>
rect -10413 25266 -10357 25268
rect -10413 25214 -10411 25266
rect -10411 25214 -10359 25266
rect -10359 25214 -10357 25266
rect -10413 25212 -10357 25214
rect -10288 25266 -10232 25268
rect -10288 25214 -10286 25266
rect -10286 25214 -10234 25266
rect -10234 25214 -10232 25266
rect -10288 25212 -10232 25214
rect -10163 25266 -10107 25268
rect -10163 25214 -10161 25266
rect -10161 25214 -10109 25266
rect -10109 25214 -10107 25266
rect -10163 25212 -10107 25214
rect -8643 25276 -8587 25278
rect -8643 25224 -8641 25276
rect -8641 25224 -8589 25276
rect -8589 25224 -8587 25276
rect -8643 25222 -8587 25224
rect -8518 25276 -8462 25278
rect -8518 25224 -8516 25276
rect -8516 25224 -8464 25276
rect -8464 25224 -8462 25276
rect -8518 25222 -8462 25224
rect -8393 25276 -8337 25278
rect -8393 25224 -8391 25276
rect -8391 25224 -8339 25276
rect -8339 25224 -8337 25276
rect -8393 25222 -8337 25224
rect -6913 25266 -6857 25268
rect -6913 25214 -6911 25266
rect -6911 25214 -6859 25266
rect -6859 25214 -6857 25266
rect -6913 25212 -6857 25214
rect -6788 25266 -6732 25268
rect -6788 25214 -6786 25266
rect -6786 25214 -6734 25266
rect -6734 25214 -6732 25266
rect -6788 25212 -6732 25214
rect -6663 25266 -6607 25268
rect -6663 25214 -6661 25266
rect -6661 25214 -6609 25266
rect -6609 25214 -6607 25266
rect -6663 25212 -6607 25214
rect -468 24621 -412 24623
rect -468 24569 -466 24621
rect -466 24569 -414 24621
rect -414 24569 -412 24621
rect -468 24567 -412 24569
rect -468 24496 -412 24498
rect -468 24444 -466 24496
rect -466 24444 -414 24496
rect -414 24444 -412 24496
rect -468 24442 -412 24444
rect -468 24371 -412 24373
rect -468 24319 -466 24371
rect -466 24319 -414 24371
rect -414 24319 -412 24371
rect -468 24317 -412 24319
rect -488 23431 -432 23433
rect -488 23379 -486 23431
rect -486 23379 -434 23431
rect -434 23379 -432 23431
rect -488 23377 -432 23379
rect -488 23306 -432 23308
rect -488 23254 -486 23306
rect -486 23254 -434 23306
rect -434 23254 -432 23306
rect -488 23252 -432 23254
rect -488 23181 -432 23183
rect -488 23129 -486 23181
rect -486 23129 -434 23181
rect -434 23129 -432 23181
rect -488 23127 -432 23129
rect 967 23266 1023 23268
rect 967 23214 969 23266
rect 969 23214 1021 23266
rect 1021 23214 1023 23266
rect 967 23212 1023 23214
rect 1092 23266 1148 23268
rect 1092 23214 1094 23266
rect 1094 23214 1146 23266
rect 1146 23214 1148 23266
rect 1092 23212 1148 23214
rect 1217 23266 1273 23268
rect 1217 23214 1219 23266
rect 1219 23214 1271 23266
rect 1271 23214 1273 23266
rect 1217 23212 1273 23214
rect 1837 23276 1893 23278
rect 1837 23224 1839 23276
rect 1839 23224 1891 23276
rect 1891 23224 1893 23276
rect 1837 23222 1893 23224
rect 1962 23276 2018 23278
rect 1962 23224 1964 23276
rect 1964 23224 2016 23276
rect 2016 23224 2018 23276
rect 1962 23222 2018 23224
rect 2087 23276 2143 23278
rect 2087 23224 2089 23276
rect 2089 23224 2141 23276
rect 2141 23224 2143 23276
rect 2087 23222 2143 23224
rect 2737 23276 2793 23278
rect 2737 23224 2739 23276
rect 2739 23224 2791 23276
rect 2791 23224 2793 23276
rect 2737 23222 2793 23224
rect 2862 23276 2918 23278
rect 2862 23224 2864 23276
rect 2864 23224 2916 23276
rect 2916 23224 2918 23276
rect 2862 23222 2918 23224
rect 2987 23276 3043 23278
rect 2987 23224 2989 23276
rect 2989 23224 3041 23276
rect 3041 23224 3043 23276
rect 2987 23222 3043 23224
rect 3637 23276 3693 23278
rect 3637 23224 3639 23276
rect 3639 23224 3691 23276
rect 3691 23224 3693 23276
rect 3637 23222 3693 23224
rect 3762 23276 3818 23278
rect 3762 23224 3764 23276
rect 3764 23224 3816 23276
rect 3816 23224 3818 23276
rect 3762 23222 3818 23224
rect 3887 23276 3943 23278
rect 3887 23224 3889 23276
rect 3889 23224 3941 23276
rect 3941 23224 3943 23276
rect 3887 23222 3943 23224
rect 4527 23276 4583 23278
rect 4527 23224 4529 23276
rect 4529 23224 4581 23276
rect 4581 23224 4583 23276
rect 4527 23222 4583 23224
rect 4652 23276 4708 23278
rect 4652 23224 4654 23276
rect 4654 23224 4706 23276
rect 4706 23224 4708 23276
rect 4652 23222 4708 23224
rect 4777 23276 4833 23278
rect 4777 23224 4779 23276
rect 4779 23224 4831 23276
rect 4831 23224 4833 23276
rect 4777 23222 4833 23224
rect 5427 23276 5483 23278
rect 5427 23224 5429 23276
rect 5429 23224 5481 23276
rect 5481 23224 5483 23276
rect 5427 23222 5483 23224
rect 5552 23276 5608 23278
rect 5552 23224 5554 23276
rect 5554 23224 5606 23276
rect 5606 23224 5608 23276
rect 5552 23222 5608 23224
rect 5677 23276 5733 23278
rect 5677 23224 5679 23276
rect 5679 23224 5731 23276
rect 5731 23224 5733 23276
rect 5677 23222 5733 23224
rect 6337 23276 6393 23278
rect 6337 23224 6339 23276
rect 6339 23224 6391 23276
rect 6391 23224 6393 23276
rect 6337 23222 6393 23224
rect 6462 23276 6518 23278
rect 6462 23224 6464 23276
rect 6464 23224 6516 23276
rect 6516 23224 6518 23276
rect 6462 23222 6518 23224
rect 6587 23276 6643 23278
rect 6587 23224 6589 23276
rect 6589 23224 6641 23276
rect 6641 23224 6643 23276
rect 6587 23222 6643 23224
rect 6967 23276 7023 23278
rect 6967 23224 6969 23276
rect 6969 23224 7021 23276
rect 7021 23224 7023 23276
rect 6967 23222 7023 23224
rect 7092 23276 7148 23278
rect 7092 23224 7094 23276
rect 7094 23224 7146 23276
rect 7146 23224 7148 23276
rect 7092 23222 7148 23224
rect 7217 23276 7273 23278
rect 7217 23224 7219 23276
rect 7219 23224 7271 23276
rect 7271 23224 7273 23276
rect 7217 23222 7273 23224
rect 8157 23276 8213 23278
rect 8157 23224 8159 23276
rect 8159 23224 8211 23276
rect 8211 23224 8213 23276
rect 8157 23222 8213 23224
rect 8282 23276 8338 23278
rect 8282 23224 8284 23276
rect 8284 23224 8336 23276
rect 8336 23224 8338 23276
rect 8282 23222 8338 23224
rect 8407 23276 8463 23278
rect 8407 23224 8409 23276
rect 8409 23224 8461 23276
rect 8461 23224 8463 23276
rect 8407 23222 8463 23224
rect 9757 23276 9813 23278
rect 9757 23224 9759 23276
rect 9759 23224 9811 23276
rect 9811 23224 9813 23276
rect 9757 23222 9813 23224
rect 9882 23276 9938 23278
rect 9882 23224 9884 23276
rect 9884 23224 9936 23276
rect 9936 23224 9938 23276
rect 9882 23222 9938 23224
rect 10007 23276 10063 23278
rect 10007 23224 10009 23276
rect 10009 23224 10061 23276
rect 10061 23224 10063 23276
rect 10007 23222 10063 23224
rect 11327 23276 11383 23278
rect 11327 23224 11329 23276
rect 11329 23224 11381 23276
rect 11381 23224 11383 23276
rect 11327 23222 11383 23224
rect 11452 23276 11508 23278
rect 11452 23224 11454 23276
rect 11454 23224 11506 23276
rect 11506 23224 11508 23276
rect 11452 23222 11508 23224
rect 11577 23276 11633 23278
rect 11577 23224 11579 23276
rect 11579 23224 11631 23276
rect 11631 23224 11633 23276
rect 11577 23222 11633 23224
rect 13047 23276 13103 23278
rect 13047 23224 13049 23276
rect 13049 23224 13101 23276
rect 13101 23224 13103 23276
rect 13047 23222 13103 23224
rect 13172 23276 13228 23278
rect 13172 23224 13174 23276
rect 13174 23224 13226 23276
rect 13226 23224 13228 23276
rect 13172 23222 13228 23224
rect 13297 23276 13353 23278
rect 13297 23224 13299 23276
rect 13299 23224 13351 23276
rect 13351 23224 13353 23276
rect 13297 23222 13353 23224
rect 15857 23266 15913 23268
rect 15857 23214 15859 23266
rect 15859 23214 15911 23266
rect 15911 23214 15913 23266
rect 15857 23212 15913 23214
rect 15982 23266 16038 23268
rect 15982 23214 15984 23266
rect 15984 23214 16036 23266
rect 16036 23214 16038 23266
rect 15982 23212 16038 23214
rect 16107 23266 16163 23268
rect 16107 23214 16109 23266
rect 16109 23214 16161 23266
rect 16161 23214 16163 23266
rect 16107 23212 16163 23214
rect 19417 23266 19473 23268
rect 19417 23214 19419 23266
rect 19419 23214 19471 23266
rect 19471 23214 19473 23266
rect 19417 23212 19473 23214
rect 19542 23266 19598 23268
rect 19542 23214 19544 23266
rect 19544 23214 19596 23266
rect 19596 23214 19598 23266
rect 19542 23212 19598 23214
rect 19667 23266 19723 23268
rect 19667 23214 19669 23266
rect 19669 23214 19721 23266
rect 19721 23214 19723 23266
rect 19667 23212 19723 23214
rect 22697 23266 22753 23268
rect 22697 23214 22699 23266
rect 22699 23214 22751 23266
rect 22751 23214 22753 23266
rect 22697 23212 22753 23214
rect 22822 23266 22878 23268
rect 22822 23214 22824 23266
rect 22824 23214 22876 23266
rect 22876 23214 22878 23266
rect 22822 23212 22878 23214
rect 22947 23266 23003 23268
rect 22947 23214 22949 23266
rect 22949 23214 23001 23266
rect 23001 23214 23003 23266
rect 22947 23212 23003 23214
rect 23242 19521 23298 19523
rect 23242 19469 23244 19521
rect 23244 19469 23296 19521
rect 23296 19469 23298 19521
rect 23242 19467 23298 19469
rect 12612 19331 12668 19333
rect 12612 19279 12614 19331
rect 12614 19279 12666 19331
rect 12666 19279 12668 19331
rect 12612 19277 12668 19279
rect 12612 19206 12668 19208
rect 12612 19154 12614 19206
rect 12614 19154 12666 19206
rect 12666 19154 12668 19206
rect 12612 19152 12668 19154
rect 23242 19396 23298 19398
rect 23242 19344 23244 19396
rect 23244 19344 23296 19396
rect 23296 19344 23298 19396
rect 23242 19342 23298 19344
rect 23242 19271 23298 19273
rect 23242 19219 23244 19271
rect 23244 19219 23296 19271
rect 23296 19219 23298 19271
rect 23242 19217 23298 19219
rect 12612 19081 12668 19083
rect 12612 19029 12614 19081
rect 12614 19029 12666 19081
rect 12666 19029 12668 19081
rect 12612 19027 12668 19029
rect 23087 18982 23143 19038
rect 12612 18601 12668 18603
rect 12612 18549 12614 18601
rect 12614 18549 12666 18601
rect 12666 18549 12668 18601
rect 12612 18547 12668 18549
rect 12612 18476 12668 18478
rect 12612 18424 12614 18476
rect 12614 18424 12666 18476
rect 12666 18424 12668 18476
rect 12612 18422 12668 18424
rect 11077 18356 11133 18358
rect 11077 18304 11079 18356
rect 11079 18304 11131 18356
rect 11131 18304 11133 18356
rect 11077 18302 11133 18304
rect 11202 18356 11258 18358
rect 11202 18304 11204 18356
rect 11204 18304 11256 18356
rect 11256 18304 11258 18356
rect 11202 18302 11258 18304
rect 12612 18351 12668 18353
rect 12612 18299 12614 18351
rect 12614 18299 12666 18351
rect 12666 18299 12668 18351
rect 12612 18297 12668 18299
rect 23712 16496 23768 16498
rect 23712 16444 23714 16496
rect 23714 16444 23766 16496
rect 23766 16444 23768 16496
rect 23712 16442 23768 16444
rect 23812 16496 23868 16498
rect 23812 16444 23814 16496
rect 23814 16444 23866 16496
rect 23866 16444 23868 16496
rect 23812 16442 23868 16444
rect 14512 16346 14568 16348
rect 14512 16294 14514 16346
rect 14514 16294 14566 16346
rect 14566 16294 14568 16346
rect 14512 16292 14568 16294
rect 14612 16346 14668 16348
rect 14612 16294 14614 16346
rect 14614 16294 14666 16346
rect 14666 16294 14668 16346
rect 14612 16292 14668 16294
rect 22312 16336 22368 16338
rect 22312 16284 22314 16336
rect 22314 16284 22366 16336
rect 22366 16284 22368 16336
rect 22312 16282 22368 16284
rect 14602 16166 14658 16168
rect 14602 16114 14604 16166
rect 14604 16114 14656 16166
rect 14656 16114 14658 16166
rect 14602 16112 14658 16114
rect 14602 16046 14658 16048
rect 14602 15994 14604 16046
rect 14604 15994 14656 16046
rect 14656 15994 14658 16046
rect 14602 15992 14658 15994
rect 15102 15906 15158 15908
rect 15102 15854 15104 15906
rect 15104 15854 15156 15906
rect 15156 15854 15158 15906
rect 15102 15852 15158 15854
rect 15102 15786 15158 15788
rect 15102 15734 15104 15786
rect 15104 15734 15156 15786
rect 15156 15734 15158 15786
rect 15102 15732 15158 15734
rect 29522 16166 29578 16168
rect 29522 16114 29524 16166
rect 29524 16114 29576 16166
rect 29576 16114 29578 16166
rect 29522 16112 29578 16114
rect 29522 16086 29578 16088
rect 29522 16034 29524 16086
rect 29524 16034 29576 16086
rect 29576 16034 29578 16086
rect 29522 16032 29578 16034
rect 29342 15906 29398 15908
rect 29342 15854 29344 15906
rect 29344 15854 29396 15906
rect 29396 15854 29398 15906
rect 29342 15852 29398 15854
rect 29342 15826 29398 15828
rect 29342 15774 29344 15826
rect 29344 15774 29396 15826
rect 29396 15774 29398 15826
rect 29342 15772 29398 15774
rect 897 14986 953 14988
rect 897 14934 899 14986
rect 899 14934 951 14986
rect 951 14934 953 14986
rect 897 14932 953 14934
rect 1022 14986 1078 14988
rect 1022 14934 1024 14986
rect 1024 14934 1076 14986
rect 1076 14934 1078 14986
rect 1022 14932 1078 14934
rect 1147 14986 1203 14988
rect 1147 14934 1149 14986
rect 1149 14934 1201 14986
rect 1201 14934 1203 14986
rect 1147 14932 1203 14934
rect 897 14866 953 14868
rect 897 14814 899 14866
rect 899 14814 951 14866
rect 951 14814 953 14866
rect 897 14812 953 14814
rect 1022 14866 1078 14868
rect 1022 14814 1024 14866
rect 1024 14814 1076 14866
rect 1076 14814 1078 14866
rect 1022 14812 1078 14814
rect 1147 14866 1203 14868
rect 1147 14814 1149 14866
rect 1149 14814 1201 14866
rect 1201 14814 1203 14866
rect 1147 14812 1203 14814
rect 2617 14986 2673 14988
rect 2617 14934 2619 14986
rect 2619 14934 2671 14986
rect 2671 14934 2673 14986
rect 2617 14932 2673 14934
rect 2742 14986 2798 14988
rect 2742 14934 2744 14986
rect 2744 14934 2796 14986
rect 2796 14934 2798 14986
rect 2742 14932 2798 14934
rect 2867 14986 2923 14988
rect 2867 14934 2869 14986
rect 2869 14934 2921 14986
rect 2921 14934 2923 14986
rect 2867 14932 2923 14934
rect 2617 14866 2673 14868
rect 2617 14814 2619 14866
rect 2619 14814 2671 14866
rect 2671 14814 2673 14866
rect 2617 14812 2673 14814
rect 2742 14866 2798 14868
rect 2742 14814 2744 14866
rect 2744 14814 2796 14866
rect 2796 14814 2798 14866
rect 2742 14812 2798 14814
rect 2867 14866 2923 14868
rect 2867 14814 2869 14866
rect 2869 14814 2921 14866
rect 2921 14814 2923 14866
rect 2867 14812 2923 14814
rect 4057 14986 4113 14988
rect 4057 14934 4059 14986
rect 4059 14934 4111 14986
rect 4111 14934 4113 14986
rect 4057 14932 4113 14934
rect 4182 14986 4238 14988
rect 4182 14934 4184 14986
rect 4184 14934 4236 14986
rect 4236 14934 4238 14986
rect 4182 14932 4238 14934
rect 4307 14986 4363 14988
rect 4307 14934 4309 14986
rect 4309 14934 4361 14986
rect 4361 14934 4363 14986
rect 4307 14932 4363 14934
rect 4057 14866 4113 14868
rect 4057 14814 4059 14866
rect 4059 14814 4111 14866
rect 4111 14814 4113 14866
rect 4057 14812 4113 14814
rect 4182 14866 4238 14868
rect 4182 14814 4184 14866
rect 4184 14814 4236 14866
rect 4236 14814 4238 14866
rect 4182 14812 4238 14814
rect 4307 14866 4363 14868
rect 4307 14814 4309 14866
rect 4309 14814 4361 14866
rect 4361 14814 4363 14866
rect 4307 14812 4363 14814
rect 5517 14986 5573 14988
rect 5517 14934 5519 14986
rect 5519 14934 5571 14986
rect 5571 14934 5573 14986
rect 5517 14932 5573 14934
rect 5642 14986 5698 14988
rect 5642 14934 5644 14986
rect 5644 14934 5696 14986
rect 5696 14934 5698 14986
rect 5642 14932 5698 14934
rect 5767 14986 5823 14988
rect 5767 14934 5769 14986
rect 5769 14934 5821 14986
rect 5821 14934 5823 14986
rect 5767 14932 5823 14934
rect 5517 14866 5573 14868
rect 5517 14814 5519 14866
rect 5519 14814 5571 14866
rect 5571 14814 5573 14866
rect 5517 14812 5573 14814
rect 5642 14866 5698 14868
rect 5642 14814 5644 14866
rect 5644 14814 5696 14866
rect 5696 14814 5698 14866
rect 5642 14812 5698 14814
rect 5767 14866 5823 14868
rect 5767 14814 5769 14866
rect 5769 14814 5821 14866
rect 5821 14814 5823 14866
rect 5767 14812 5823 14814
rect 7357 14946 7413 14948
rect 7357 14894 7359 14946
rect 7359 14894 7411 14946
rect 7411 14894 7413 14946
rect 7357 14892 7413 14894
rect 7482 14946 7538 14948
rect 7482 14894 7484 14946
rect 7484 14894 7536 14946
rect 7536 14894 7538 14946
rect 7482 14892 7538 14894
rect 7607 14946 7663 14948
rect 7607 14894 7609 14946
rect 7609 14894 7661 14946
rect 7661 14894 7663 14946
rect 7607 14892 7663 14894
rect 8827 14956 8883 14958
rect 8827 14904 8829 14956
rect 8829 14904 8881 14956
rect 8881 14904 8883 14956
rect 8827 14902 8883 14904
rect 8952 14956 9008 14958
rect 8952 14904 8954 14956
rect 8954 14904 9006 14956
rect 9006 14904 9008 14956
rect 8952 14902 9008 14904
rect 9077 14956 9133 14958
rect 9077 14904 9079 14956
rect 9079 14904 9131 14956
rect 9131 14904 9133 14956
rect 9077 14902 9133 14904
rect 11687 14966 11743 14968
rect 11687 14914 11689 14966
rect 11689 14914 11741 14966
rect 11741 14914 11743 14966
rect 11687 14912 11743 14914
rect 11812 14966 11868 14968
rect 11812 14914 11814 14966
rect 11814 14914 11866 14966
rect 11866 14914 11868 14966
rect 11812 14912 11868 14914
rect 11937 14966 11993 14968
rect 11937 14914 11939 14966
rect 11939 14914 11991 14966
rect 11991 14914 11993 14966
rect 11937 14912 11993 14914
rect 12697 14966 12753 14968
rect 12697 14914 12699 14966
rect 12699 14914 12751 14966
rect 12751 14914 12753 14966
rect 12697 14912 12753 14914
rect 12822 14966 12878 14968
rect 12822 14914 12824 14966
rect 12824 14914 12876 14966
rect 12876 14914 12878 14966
rect 12822 14912 12878 14914
rect 12947 14966 13003 14968
rect 12947 14914 12949 14966
rect 12949 14914 13001 14966
rect 13001 14914 13003 14966
rect 12947 14912 13003 14914
rect 14602 14956 14658 14958
rect 14602 14904 14604 14956
rect 14604 14904 14656 14956
rect 14656 14904 14658 14956
rect 14602 14902 14658 14904
rect 15267 14966 15323 14968
rect 15267 14914 15269 14966
rect 15269 14914 15321 14966
rect 15321 14914 15323 14966
rect 15267 14912 15323 14914
rect 15392 14966 15448 14968
rect 15392 14914 15394 14966
rect 15394 14914 15446 14966
rect 15446 14914 15448 14966
rect 15392 14912 15448 14914
rect 15517 14966 15573 14968
rect 15517 14914 15519 14966
rect 15519 14914 15571 14966
rect 15571 14914 15573 14966
rect 15517 14912 15573 14914
rect 15747 14966 15803 14968
rect 15747 14914 15749 14966
rect 15749 14914 15801 14966
rect 15801 14914 15803 14966
rect 15747 14912 15803 14914
rect 15872 14966 15928 14968
rect 15872 14914 15874 14966
rect 15874 14914 15926 14966
rect 15926 14914 15928 14966
rect 15872 14912 15928 14914
rect 15997 14966 16053 14968
rect 15997 14914 15999 14966
rect 15999 14914 16051 14966
rect 16051 14914 16053 14966
rect 15997 14912 16053 14914
rect 20527 14946 20583 14948
rect 20527 14894 20529 14946
rect 20529 14894 20581 14946
rect 20581 14894 20583 14946
rect 20527 14892 20583 14894
rect 20652 14946 20708 14948
rect 20652 14894 20654 14946
rect 20654 14894 20706 14946
rect 20706 14894 20708 14946
rect 20652 14892 20708 14894
rect 20777 14946 20833 14948
rect 20777 14894 20779 14946
rect 20779 14894 20831 14946
rect 20831 14894 20833 14946
rect 20777 14892 20833 14894
rect 20887 14946 20943 14948
rect 20887 14894 20889 14946
rect 20889 14894 20941 14946
rect 20941 14894 20943 14946
rect 20887 14892 20943 14894
rect 21012 14946 21068 14948
rect 21012 14894 21014 14946
rect 21014 14894 21066 14946
rect 21066 14894 21068 14946
rect 21012 14892 21068 14894
rect 21137 14946 21193 14948
rect 21137 14894 21139 14946
rect 21139 14894 21191 14946
rect 21191 14894 21193 14946
rect 21137 14892 21193 14894
rect 16092 14472 16148 14528
rect 20272 14526 20328 14528
rect 20272 14474 20274 14526
rect 20274 14474 20326 14526
rect 20326 14474 20328 14526
rect 20272 14472 20328 14474
rect 22312 14196 22368 14198
rect 22312 14144 22314 14196
rect 22314 14144 22366 14196
rect 22366 14144 22368 14196
rect 22312 14142 22368 14144
rect 21252 14002 21308 14058
rect -6978 12906 -6922 12908
rect -6978 12854 -6976 12906
rect -6976 12854 -6924 12906
rect -6924 12854 -6922 12906
rect -6978 12852 -6922 12854
rect -7348 12766 -7292 12768
rect -7348 12714 -7346 12766
rect -7346 12714 -7294 12766
rect -7294 12714 -7292 12766
rect -7348 12712 -7292 12714
rect -10878 12642 -10822 12698
rect -10738 12532 -10682 12588
rect -10458 12342 -10402 12398
rect -10318 12232 -10262 12288
rect -6148 12047 -6092 12103
rect -6058 12047 -6002 12103
rect -6358 11807 -6302 11863
rect -6268 11807 -6212 11863
rect -6578 11456 -6522 11458
rect -6578 11404 -6576 11456
rect -6576 11404 -6524 11456
rect -6524 11404 -6522 11456
rect -6578 11402 -6522 11404
rect -6458 11456 -6402 11458
rect -6458 11404 -6456 11456
rect -6456 11404 -6404 11456
rect -6404 11404 -6402 11456
rect -6458 11402 -6402 11404
rect 957 7476 1013 7478
rect 957 7424 959 7476
rect 959 7424 1011 7476
rect 1011 7424 1013 7476
rect 957 7422 1013 7424
rect 1082 7476 1138 7478
rect 1082 7424 1084 7476
rect 1084 7424 1136 7476
rect 1136 7424 1138 7476
rect 1082 7422 1138 7424
rect 1567 7476 1623 7478
rect 1567 7424 1569 7476
rect 1569 7424 1621 7476
rect 1621 7424 1623 7476
rect 1567 7422 1623 7424
rect 1692 7476 1748 7478
rect 1692 7424 1694 7476
rect 1694 7424 1746 7476
rect 1746 7424 1748 7476
rect 1692 7422 1748 7424
rect 2717 7476 2773 7478
rect 2717 7424 2719 7476
rect 2719 7424 2771 7476
rect 2771 7424 2773 7476
rect 2717 7422 2773 7424
rect 2842 7476 2898 7478
rect 2842 7424 2844 7476
rect 2844 7424 2896 7476
rect 2896 7424 2898 7476
rect 2842 7422 2898 7424
rect 3887 7476 3943 7478
rect 3887 7424 3889 7476
rect 3889 7424 3941 7476
rect 3941 7424 3943 7476
rect 3887 7422 3943 7424
rect 4012 7476 4068 7478
rect 4012 7424 4014 7476
rect 4014 7424 4066 7476
rect 4066 7424 4068 7476
rect 4012 7422 4068 7424
rect 5047 7476 5103 7478
rect 5047 7424 5049 7476
rect 5049 7424 5101 7476
rect 5101 7424 5103 7476
rect 5047 7422 5103 7424
rect 5172 7476 5228 7478
rect 5172 7424 5174 7476
rect 5174 7424 5226 7476
rect 5226 7424 5228 7476
rect 5172 7422 5228 7424
rect 6217 7476 6273 7478
rect 6217 7424 6219 7476
rect 6219 7424 6271 7476
rect 6271 7424 6273 7476
rect 6217 7422 6273 7424
rect 6342 7476 6398 7478
rect 6342 7424 6344 7476
rect 6344 7424 6396 7476
rect 6396 7424 6398 7476
rect 6342 7422 6398 7424
rect 7377 7476 7433 7478
rect 7377 7424 7379 7476
rect 7379 7424 7431 7476
rect 7431 7424 7433 7476
rect 7377 7422 7433 7424
rect 7502 7476 7558 7478
rect 7502 7424 7504 7476
rect 7504 7424 7556 7476
rect 7556 7424 7558 7476
rect 7502 7422 7558 7424
rect 1397 406 1453 408
rect 1397 354 1399 406
rect 1399 354 1451 406
rect 1451 354 1453 406
rect 1397 352 1453 354
rect 1522 406 1578 408
rect 1522 354 1524 406
rect 1524 354 1576 406
rect 1576 354 1578 406
rect 1522 352 1578 354
rect 1647 406 1703 408
rect 1647 354 1649 406
rect 1649 354 1701 406
rect 1701 354 1703 406
rect 1647 352 1703 354
rect 3127 406 3183 408
rect 3127 354 3129 406
rect 3129 354 3181 406
rect 3181 354 3183 406
rect 3127 352 3183 354
rect 3252 406 3308 408
rect 3252 354 3254 406
rect 3254 354 3306 406
rect 3306 354 3308 406
rect 3252 352 3308 354
rect 3377 406 3433 408
rect 3377 354 3379 406
rect 3379 354 3431 406
rect 3431 354 3433 406
rect 3377 352 3433 354
rect 5187 406 5243 408
rect 5187 354 5189 406
rect 5189 354 5241 406
rect 5241 354 5243 406
rect 5187 352 5243 354
rect 5312 406 5368 408
rect 5312 354 5314 406
rect 5314 354 5366 406
rect 5366 354 5368 406
rect 5312 352 5368 354
rect 5437 406 5493 408
rect 5437 354 5439 406
rect 5439 354 5491 406
rect 5491 354 5493 406
rect 5437 352 5493 354
rect 8827 396 8883 398
rect 8827 344 8829 396
rect 8829 344 8881 396
rect 8881 344 8883 396
rect 8827 342 8883 344
rect 8952 396 9008 398
rect 8952 344 8954 396
rect 8954 344 9006 396
rect 9006 344 9008 396
rect 8952 342 9008 344
rect 9077 396 9133 398
rect 9077 344 9079 396
rect 9079 344 9131 396
rect 9131 344 9133 396
rect 9077 342 9133 344
rect 10947 396 11003 398
rect 10947 344 10949 396
rect 10949 344 11001 396
rect 11001 344 11003 396
rect 10947 342 11003 344
rect 11072 396 11128 398
rect 11072 344 11074 396
rect 11074 344 11126 396
rect 11126 344 11128 396
rect 11072 342 11128 344
rect 11197 396 11253 398
rect 11197 344 11199 396
rect 11199 344 11251 396
rect 11251 344 11253 396
rect 11197 342 11253 344
rect 14677 396 14733 398
rect 14677 344 14679 396
rect 14679 344 14731 396
rect 14731 344 14733 396
rect 14677 342 14733 344
rect 14802 396 14858 398
rect 14802 344 14804 396
rect 14804 344 14856 396
rect 14856 344 14858 396
rect 14802 342 14858 344
rect 14927 396 14983 398
rect 14927 344 14929 396
rect 14929 344 14981 396
rect 14981 344 14983 396
rect 14927 342 14983 344
rect 17037 396 17093 398
rect 17037 344 17039 396
rect 17039 344 17091 396
rect 17091 344 17093 396
rect 17037 342 17093 344
rect 17162 396 17218 398
rect 17162 344 17164 396
rect 17164 344 17216 396
rect 17216 344 17218 396
rect 17162 342 17218 344
rect 17287 396 17343 398
rect 17287 344 17289 396
rect 17289 344 17341 396
rect 17341 344 17343 396
rect 17287 342 17343 344
rect 19047 396 19103 398
rect 19047 344 19049 396
rect 19049 344 19101 396
rect 19101 344 19103 396
rect 19047 342 19103 344
rect 19172 396 19228 398
rect 19172 344 19174 396
rect 19174 344 19226 396
rect 19226 344 19228 396
rect 19172 342 19228 344
rect 19297 396 19353 398
rect 19297 344 19299 396
rect 19299 344 19351 396
rect 19351 344 19353 396
rect 19297 342 19353 344
rect 21007 396 21063 398
rect 21007 344 21009 396
rect 21009 344 21061 396
rect 21061 344 21063 396
rect 21007 342 21063 344
rect 21132 396 21188 398
rect 21132 344 21134 396
rect 21134 344 21186 396
rect 21186 344 21188 396
rect 21132 342 21188 344
rect 21257 396 21313 398
rect 21257 344 21259 396
rect 21259 344 21311 396
rect 21311 344 21313 396
rect 21257 342 21313 344
<< metal3 >>
rect -10440 25272 -10080 25300
rect -10440 25208 -10417 25272
rect -10353 25208 -10292 25272
rect -10228 25208 -10167 25272
rect -10103 25208 -10080 25272
rect -10440 25180 -10080 25208
rect -8670 25282 -8310 25310
rect -8670 25218 -8647 25282
rect -8583 25218 -8522 25282
rect -8458 25218 -8397 25282
rect -8333 25218 -8310 25282
rect -8670 25190 -8310 25218
rect -6940 25272 -6580 25300
rect -6940 25208 -6917 25272
rect -6853 25208 -6792 25272
rect -6728 25208 -6667 25272
rect -6603 25208 -6580 25272
rect -6940 25180 -6580 25208
rect -500 24627 -380 24650
rect -500 24563 -472 24627
rect -408 24563 -380 24627
rect -500 24502 -380 24563
rect -500 24438 -472 24502
rect -408 24438 -380 24502
rect -500 24377 -380 24438
rect -500 24313 -472 24377
rect -408 24313 -380 24377
rect -500 24290 -380 24313
rect -520 23437 -400 23460
rect -520 23373 -492 23437
rect -428 23373 -400 23437
rect -520 23312 -400 23373
rect -520 23248 -492 23312
rect -428 23248 -400 23312
rect -520 23187 -400 23248
rect -520 23123 -492 23187
rect -428 23123 -400 23187
rect 940 23272 1300 23300
rect 940 23208 963 23272
rect 1027 23208 1088 23272
rect 1152 23208 1213 23272
rect 1277 23208 1300 23272
rect 940 23180 1300 23208
rect 1810 23282 2170 23310
rect 1810 23218 1833 23282
rect 1897 23218 1958 23282
rect 2022 23218 2083 23282
rect 2147 23218 2170 23282
rect 1810 23190 2170 23218
rect 2710 23282 3070 23310
rect 2710 23218 2733 23282
rect 2797 23218 2858 23282
rect 2922 23218 2983 23282
rect 3047 23218 3070 23282
rect 2710 23190 3070 23218
rect 3610 23282 3970 23310
rect 3610 23218 3633 23282
rect 3697 23218 3758 23282
rect 3822 23218 3883 23282
rect 3947 23218 3970 23282
rect 3610 23190 3970 23218
rect 4500 23282 4860 23310
rect 4500 23218 4523 23282
rect 4587 23218 4648 23282
rect 4712 23218 4773 23282
rect 4837 23218 4860 23282
rect 4500 23190 4860 23218
rect 5400 23282 5760 23310
rect 5400 23218 5423 23282
rect 5487 23218 5548 23282
rect 5612 23218 5673 23282
rect 5737 23218 5760 23282
rect 5400 23190 5760 23218
rect 6310 23282 6670 23310
rect 6310 23218 6333 23282
rect 6397 23218 6458 23282
rect 6522 23218 6583 23282
rect 6647 23218 6670 23282
rect 6310 23190 6670 23218
rect 6940 23282 7300 23310
rect 6940 23218 6963 23282
rect 7027 23218 7088 23282
rect 7152 23218 7213 23282
rect 7277 23218 7300 23282
rect 6940 23190 7300 23218
rect 8130 23282 8490 23310
rect 8130 23218 8153 23282
rect 8217 23218 8278 23282
rect 8342 23218 8403 23282
rect 8467 23218 8490 23282
rect 8130 23190 8490 23218
rect 9730 23282 10090 23310
rect 9730 23218 9753 23282
rect 9817 23218 9878 23282
rect 9942 23218 10003 23282
rect 10067 23218 10090 23282
rect 9730 23190 10090 23218
rect 11300 23282 11660 23310
rect 11300 23218 11323 23282
rect 11387 23218 11448 23282
rect 11512 23218 11573 23282
rect 11637 23218 11660 23282
rect 11300 23190 11660 23218
rect 13020 23282 13380 23310
rect 13020 23218 13043 23282
rect 13107 23218 13168 23282
rect 13232 23218 13293 23282
rect 13357 23218 13380 23282
rect 13020 23190 13380 23218
rect 15830 23272 16190 23300
rect 15830 23208 15853 23272
rect 15917 23208 15978 23272
rect 16042 23208 16103 23272
rect 16167 23208 16190 23272
rect 15830 23180 16190 23208
rect 19390 23272 19750 23300
rect 19390 23208 19413 23272
rect 19477 23208 19538 23272
rect 19602 23208 19663 23272
rect 19727 23208 19750 23272
rect 19390 23180 19750 23208
rect 22670 23272 23030 23300
rect 22670 23208 22693 23272
rect 22757 23208 22818 23272
rect 22882 23208 22943 23272
rect 23007 23208 23030 23272
rect 22670 23180 23030 23208
rect -520 23100 -400 23123
rect -10890 12698 -10810 20840
rect -10890 12642 -10878 12698
rect -10822 12642 -10810 12698
rect -10890 12630 -10810 12642
rect -10750 12588 -10670 20800
rect -10610 12782 -10530 20820
rect -10610 12718 -10607 12782
rect -10543 12718 -10530 12782
rect -10610 12700 -10530 12718
rect -10750 12532 -10738 12588
rect -10682 12532 -10670 12588
rect -10750 12520 -10670 12532
rect -10470 12398 -10390 20800
rect -10470 12342 -10458 12398
rect -10402 12342 -10390 12398
rect -10470 12330 -10390 12342
rect -10330 12288 -10250 20800
rect 23210 19527 23330 19550
rect 23210 19463 23238 19527
rect 23302 19463 23330 19527
rect 23210 19402 23330 19463
rect 12580 19337 12700 19360
rect 12580 19273 12608 19337
rect 12672 19273 12700 19337
rect 12580 19212 12700 19273
rect 12580 19148 12608 19212
rect 12672 19148 12700 19212
rect 23210 19338 23238 19402
rect 23302 19338 23330 19402
rect 23210 19277 23330 19338
rect 23210 19213 23238 19277
rect 23302 19213 23330 19277
rect 23210 19190 23330 19213
rect 12580 19087 12700 19148
rect 12580 19023 12608 19087
rect 12672 19023 12700 19087
rect 12580 19000 12700 19023
rect 23070 19038 23160 19060
rect 23070 18982 23087 19038
rect 23143 18982 23160 19038
rect 23070 18960 23160 18982
rect 17920 18750 18270 18830
rect 12580 18607 12700 18630
rect 12580 18543 12608 18607
rect 12672 18543 12700 18607
rect 12580 18482 12700 18543
rect 12580 18418 12608 18482
rect 12672 18418 12700 18482
rect 11050 18362 11290 18390
rect 11050 18298 11073 18362
rect 11137 18298 11198 18362
rect 11262 18298 11290 18362
rect 11050 18270 11290 18298
rect 12580 18357 12700 18418
rect 12580 18293 12608 18357
rect 12672 18293 12700 18357
rect 12580 18270 12700 18293
rect 12480 18092 12610 18110
rect 12480 18028 12513 18092
rect 12577 18028 12610 18092
rect 12480 17262 12610 18028
rect 23440 17960 23680 18060
rect 12480 17198 12513 17262
rect 12577 17198 12610 17262
rect 12480 15702 12610 17198
rect 12480 15638 12513 15702
rect 12577 15638 12610 15702
rect 12480 15512 12610 15638
rect 12480 15448 12513 15512
rect 12577 15448 12610 15512
rect 12480 15420 12610 15448
rect 12670 17672 12800 17690
rect 12670 17608 12703 17672
rect 12767 17608 12800 17672
rect 12670 15320 12800 17608
rect 23580 16520 23680 17960
rect 23580 16498 23890 16520
rect 23580 16442 23712 16498
rect 23768 16442 23812 16498
rect 23868 16442 23890 16498
rect 23580 16420 23890 16442
rect 14500 16348 14680 16360
rect 14500 16292 14512 16348
rect 14568 16292 14612 16348
rect 14668 16292 14680 16348
rect 14500 16280 14680 16292
rect 22280 16338 22400 16420
rect 22280 16282 22312 16338
rect 22368 16282 22400 16338
rect 22280 16270 22400 16282
rect 14580 16172 14680 16190
rect 14580 16108 14598 16172
rect 14662 16108 14680 16172
rect 14580 16052 14680 16108
rect 14580 15988 14598 16052
rect 14662 15988 14680 16052
rect 23830 16132 24050 16190
rect 23830 16068 23848 16132
rect 23912 16068 23968 16132
rect 24032 16068 24050 16132
rect 23830 16010 24050 16068
rect 29500 16168 29600 16190
rect 29500 16132 29522 16168
rect 29578 16132 29600 16168
rect 29500 16068 29518 16132
rect 29582 16068 29600 16132
rect 29500 16032 29522 16068
rect 29578 16032 29600 16068
rect 29500 16010 29600 16032
rect 14580 15970 14680 15988
rect 15080 15912 15180 15930
rect 15080 15848 15098 15912
rect 15162 15848 15180 15912
rect 15080 15792 15180 15848
rect 15080 15728 15098 15792
rect 15162 15728 15180 15792
rect 15080 15710 15180 15728
rect 12560 15302 12800 15320
rect 12560 15238 12583 15302
rect 12647 15238 12713 15302
rect 12777 15238 12800 15302
rect 12560 15222 12800 15238
rect 12560 15158 12583 15222
rect 12647 15158 12713 15222
rect 12777 15158 12800 15222
rect 12560 15140 12800 15158
rect -490 15052 -190 15080
rect -490 14988 -462 15052
rect -398 14988 -282 15052
rect -218 14988 -190 15052
rect -490 14872 -190 14988
rect -490 14808 -462 14872
rect -398 14808 -282 14872
rect -218 14808 -190 14872
rect -7000 12912 -6900 12930
rect -7000 12848 -6982 12912
rect -6918 12848 -6900 12912
rect -7000 12830 -6900 12848
rect -7370 12772 -7270 12790
rect -7370 12708 -7352 12772
rect -7288 12708 -7270 12772
rect -7370 12690 -7270 12708
rect -10330 12232 -10318 12288
rect -10262 12232 -10250 12288
rect -10330 12220 -10250 12232
rect -5430 12542 -5190 12570
rect -5430 12478 -5402 12542
rect -5338 12478 -5282 12542
rect -5218 12478 -5190 12542
rect -5430 12450 -5190 12478
rect -6170 12103 -5990 12120
rect -6170 12047 -6148 12103
rect -6092 12047 -6058 12103
rect -6002 12047 -5990 12103
rect -6170 12020 -5990 12047
rect -6380 11863 -6190 11880
rect -6380 11807 -6358 11863
rect -6302 11807 -6268 11863
rect -6212 11807 -6190 11863
rect -6380 11780 -6190 11807
rect -6600 11462 -6380 11480
rect -6600 11398 -6582 11462
rect -6518 11398 -6462 11462
rect -6398 11398 -6380 11462
rect -6600 11380 -6380 11398
rect -7330 11222 -7110 11250
rect -7330 11158 -7312 11222
rect -7248 11158 -7192 11222
rect -7128 11158 -7110 11222
rect -7330 11130 -7110 11158
rect -6290 1140 -6190 11780
rect -6520 1040 -6190 1140
rect -6090 1040 -5990 12020
rect -5850 11042 -5610 11070
rect -5850 10978 -5822 11042
rect -5758 10978 -5702 11042
rect -5638 10978 -5610 11042
rect -5850 10950 -5610 10978
rect -5730 9020 -5610 10950
rect -5430 10520 -5310 12450
rect -5250 12362 -5010 12390
rect -5250 12298 -5222 12362
rect -5158 12298 -5102 12362
rect -5038 12298 -5010 12362
rect -5250 12270 -5010 12298
rect -5250 10862 -5130 12270
rect -5250 10798 -5222 10862
rect -5158 10798 -5130 10862
rect -5250 10770 -5130 10798
rect -5070 12172 -4830 12200
rect -5070 12108 -5042 12172
rect -4978 12108 -4922 12172
rect -4858 12108 -4830 12172
rect -5070 12080 -4830 12108
rect -5070 10700 -4950 12080
rect -5190 10672 -4950 10700
rect -5190 10608 -5162 10672
rect -5098 10608 -5042 10672
rect -4978 10608 -4950 10672
rect -5190 10580 -4950 10608
rect -490 11462 -190 14808
rect 870 14992 1230 15020
rect 870 14928 893 14992
rect 957 14928 1018 14992
rect 1082 14928 1143 14992
rect 1207 14928 1230 14992
rect 870 14872 1230 14928
rect 870 14808 893 14872
rect 957 14808 1018 14872
rect 1082 14808 1143 14872
rect 1207 14808 1230 14872
rect 870 14780 1230 14808
rect 2590 14992 2950 15020
rect 2590 14928 2613 14992
rect 2677 14928 2738 14992
rect 2802 14928 2863 14992
rect 2927 14928 2950 14992
rect 2590 14872 2950 14928
rect 2590 14808 2613 14872
rect 2677 14808 2738 14872
rect 2802 14808 2863 14872
rect 2927 14808 2950 14872
rect 2590 14780 2950 14808
rect 4030 14992 4390 15020
rect 4030 14928 4053 14992
rect 4117 14928 4178 14992
rect 4242 14928 4303 14992
rect 4367 14928 4390 14992
rect 4030 14872 4390 14928
rect 4030 14808 4053 14872
rect 4117 14808 4178 14872
rect 4242 14808 4303 14872
rect 4367 14808 4390 14872
rect 4030 14780 4390 14808
rect 5490 14992 5850 15020
rect 5490 14928 5513 14992
rect 5577 14928 5638 14992
rect 5702 14928 5763 14992
rect 5827 14928 5850 14992
rect 5490 14872 5850 14928
rect 5490 14808 5513 14872
rect 5577 14808 5638 14872
rect 5702 14808 5763 14872
rect 5827 14808 5850 14872
rect 7330 14952 7690 14980
rect 7330 14888 7353 14952
rect 7417 14888 7478 14952
rect 7542 14888 7603 14952
rect 7667 14888 7690 14952
rect 7330 14860 7690 14888
rect 8800 14962 9160 14990
rect 8800 14898 8823 14962
rect 8887 14898 8948 14962
rect 9012 14898 9073 14962
rect 9137 14898 9160 14962
rect 8800 14870 9160 14898
rect 11660 14972 12020 15000
rect 11660 14908 11683 14972
rect 11747 14908 11808 14972
rect 11872 14908 11933 14972
rect 11997 14908 12020 14972
rect 11660 14880 12020 14908
rect 12670 14972 13030 15000
rect 12670 14908 12693 14972
rect 12757 14908 12818 14972
rect 12882 14908 12943 14972
rect 13007 14908 13030 14972
rect 15240 14972 15600 15000
rect 12670 14880 13030 14908
rect 14580 14958 14680 14970
rect 14580 14902 14602 14958
rect 14658 14902 14680 14958
rect 14580 14890 14680 14902
rect 15240 14908 15263 14972
rect 15327 14908 15388 14972
rect 15452 14908 15513 14972
rect 15577 14908 15600 14972
rect 15240 14880 15600 14908
rect 15720 14972 16080 15000
rect 15720 14908 15743 14972
rect 15807 14908 15868 14972
rect 15932 14908 15993 14972
rect 16057 14908 16080 14972
rect 15720 14880 16080 14908
rect 20500 14952 21220 14980
rect 20500 14888 20523 14952
rect 20587 14888 20648 14952
rect 20712 14888 20773 14952
rect 20837 14888 20883 14952
rect 20947 14888 21008 14952
rect 21072 14888 21133 14952
rect 21197 14888 21220 14952
rect 20500 14860 21220 14888
rect 5490 14780 5850 14808
rect 16070 14532 16170 14550
rect 16070 14468 16088 14532
rect 16152 14468 16170 14532
rect 16070 14450 16170 14468
rect 20250 14532 20350 14550
rect 20250 14468 20268 14532
rect 20332 14468 20350 14532
rect 20250 14450 20350 14468
rect 21240 14058 21320 14430
rect 23950 14382 24050 16010
rect 23950 14318 23968 14382
rect 24032 14318 24050 14382
rect 23950 14262 24050 14318
rect 22280 14202 22400 14220
rect 22280 14138 22308 14202
rect 22372 14138 22400 14202
rect 23950 14198 23968 14262
rect 24032 14198 24050 14262
rect 23950 14180 24050 14198
rect 24150 15872 24370 15930
rect 24150 15808 24168 15872
rect 24232 15808 24288 15872
rect 24352 15808 24370 15872
rect 24150 15750 24370 15808
rect 29320 15908 29420 15930
rect 29320 15872 29342 15908
rect 29398 15872 29420 15908
rect 29320 15808 29338 15872
rect 29402 15808 29420 15872
rect 29320 15772 29342 15808
rect 29398 15772 29420 15808
rect 29320 15750 29420 15772
rect 24150 14382 24250 15750
rect 26750 15542 26940 15600
rect 26750 15478 26763 15542
rect 26827 15478 26863 15542
rect 26927 15478 26940 15542
rect 26750 15420 26940 15478
rect 26510 15262 26701 15320
rect 26510 15198 26523 15262
rect 26587 15198 26623 15262
rect 26687 15198 26701 15262
rect 26510 15140 26701 15198
rect 24150 14318 24168 14382
rect 24232 14318 24250 14382
rect 24150 14262 24250 14318
rect 24150 14198 24168 14262
rect 24232 14198 24250 14262
rect 24150 14180 24250 14198
rect 26599 14180 26701 15140
rect 26810 14377 26910 15420
rect 26810 14313 26828 14377
rect 26892 14313 26910 14377
rect 26810 14300 26910 14313
rect 22280 14120 22400 14138
rect 21240 14002 21252 14058
rect 21308 14002 21320 14058
rect 21240 13990 21320 14002
rect 230 13842 470 13870
rect 230 13778 258 13842
rect 322 13778 378 13842
rect 442 13778 470 13842
rect 230 13750 470 13778
rect 230 12570 350 13750
rect 110 12542 350 12570
rect 110 12478 138 12542
rect 202 12478 258 12542
rect 322 12478 350 12542
rect 110 12450 350 12478
rect 410 13662 650 13690
rect 410 13598 438 13662
rect 502 13598 558 13662
rect 622 13598 650 13662
rect 410 13570 650 13598
rect 410 12390 530 13570
rect 290 12362 530 12390
rect 290 12298 318 12362
rect 382 12298 438 12362
rect 502 12298 530 12362
rect 290 12270 530 12298
rect 590 13472 830 13500
rect 590 13408 618 13472
rect 682 13408 738 13472
rect 802 13408 830 13472
rect 590 13380 830 13408
rect 590 12200 710 13380
rect 470 12172 710 12200
rect 470 12108 498 12172
rect 562 12108 618 12172
rect 682 12108 710 12172
rect 470 12080 710 12108
rect -490 11398 -442 11462
rect -378 11398 -312 11462
rect -248 11398 -190 11462
rect -5550 10492 -5310 10520
rect -5550 10428 -5522 10492
rect -5458 10428 -5402 10492
rect -5338 10428 -5310 10492
rect -5550 10400 -5310 10428
rect -5730 8992 -5490 9020
rect -5730 8928 -5707 8992
rect -5643 8928 -5577 8992
rect -5513 8928 -5490 8992
rect -5730 8900 -5490 8928
rect -490 7572 -190 11398
rect 240 8992 480 9020
rect 240 8928 263 8992
rect 327 8928 393 8992
rect 457 8928 480 8992
rect 240 8900 480 8928
rect -490 7508 -462 7572
rect -398 7508 -282 7572
rect -218 7508 -190 7572
rect -490 7392 -190 7508
rect -490 7328 -462 7392
rect -398 7328 -282 7392
rect -218 7328 -190 7392
rect -6590 987 -6350 1040
rect -6590 923 -6567 987
rect -6503 923 -6447 987
rect -6383 923 -6350 987
rect -6590 870 -6350 923
rect -6110 977 -5860 1040
rect -6110 913 -6077 977
rect -6013 913 -5947 977
rect -5883 913 -5860 977
rect -6110 870 -5860 913
rect -6090 860 -5990 870
rect -490 472 -190 7328
rect 360 6830 480 8900
rect 930 7482 1170 7510
rect 930 7418 953 7482
rect 1017 7418 1078 7482
rect 1142 7418 1170 7482
rect 930 7390 1170 7418
rect 1540 7482 1780 7510
rect 1540 7418 1563 7482
rect 1627 7418 1688 7482
rect 1752 7418 1780 7482
rect 1540 7390 1780 7418
rect 2690 7482 2930 7510
rect 2690 7418 2713 7482
rect 2777 7418 2838 7482
rect 2902 7418 2930 7482
rect 2690 7390 2930 7418
rect 3860 7482 4100 7510
rect 3860 7418 3883 7482
rect 3947 7418 4008 7482
rect 4072 7418 4100 7482
rect 3860 7390 4100 7418
rect 5020 7482 5260 7510
rect 5020 7418 5043 7482
rect 5107 7418 5168 7482
rect 5232 7418 5260 7482
rect 5020 7390 5260 7418
rect 6190 7482 6430 7510
rect 6190 7418 6213 7482
rect 6277 7418 6338 7482
rect 6402 7418 6430 7482
rect 6190 7390 6430 7418
rect 7350 7482 7590 7510
rect 7350 7418 7373 7482
rect 7437 7418 7498 7482
rect 7562 7418 7590 7482
rect 7350 7390 7590 7418
rect 360 6812 560 6830
rect 360 6748 373 6812
rect 437 6748 483 6812
rect 547 6748 560 6812
rect 360 6730 560 6748
rect 22290 3957 22390 3970
rect 22290 3893 22308 3957
rect 22372 3893 22390 3957
rect 22290 3880 22390 3893
rect -490 408 -462 472
rect -398 408 -282 472
rect -218 408 -190 472
rect -490 292 -190 408
rect 1370 412 1730 440
rect 1370 348 1393 412
rect 1457 348 1518 412
rect 1582 348 1643 412
rect 1707 348 1730 412
rect 1370 320 1730 348
rect 3100 412 3460 440
rect 3100 348 3123 412
rect 3187 348 3248 412
rect 3312 348 3373 412
rect 3437 348 3460 412
rect 3100 320 3460 348
rect 5160 412 5520 440
rect 5160 348 5183 412
rect 5247 348 5308 412
rect 5372 348 5433 412
rect 5497 348 5520 412
rect 5160 320 5520 348
rect 8800 402 9160 430
rect 8800 338 8823 402
rect 8887 338 8948 402
rect 9012 338 9073 402
rect 9137 338 9160 402
rect 8800 310 9160 338
rect 10920 402 11280 430
rect 10920 338 10943 402
rect 11007 338 11068 402
rect 11132 338 11193 402
rect 11257 338 11280 402
rect 10920 310 11280 338
rect 14650 402 15010 430
rect 14650 338 14673 402
rect 14737 338 14798 402
rect 14862 338 14923 402
rect 14987 338 15010 402
rect 14650 310 15010 338
rect 17010 402 17370 430
rect 17010 338 17033 402
rect 17097 338 17158 402
rect 17222 338 17283 402
rect 17347 338 17370 402
rect 17010 310 17370 338
rect 19020 402 19380 430
rect 19020 338 19043 402
rect 19107 338 19168 402
rect 19232 338 19293 402
rect 19357 338 19380 402
rect 19020 310 19380 338
rect 20980 402 21340 430
rect 20980 338 21003 402
rect 21067 338 21128 402
rect 21192 338 21253 402
rect 21317 338 21340 402
rect 20980 310 21340 338
rect -490 228 -462 292
rect -398 228 -282 292
rect -218 228 -190 292
rect -490 200 -190 228
<< via3 >>
rect -10417 25268 -10353 25272
rect -10417 25212 -10413 25268
rect -10413 25212 -10357 25268
rect -10357 25212 -10353 25268
rect -10417 25208 -10353 25212
rect -10292 25268 -10228 25272
rect -10292 25212 -10288 25268
rect -10288 25212 -10232 25268
rect -10232 25212 -10228 25268
rect -10292 25208 -10228 25212
rect -10167 25268 -10103 25272
rect -10167 25212 -10163 25268
rect -10163 25212 -10107 25268
rect -10107 25212 -10103 25268
rect -10167 25208 -10103 25212
rect -8647 25278 -8583 25282
rect -8647 25222 -8643 25278
rect -8643 25222 -8587 25278
rect -8587 25222 -8583 25278
rect -8647 25218 -8583 25222
rect -8522 25278 -8458 25282
rect -8522 25222 -8518 25278
rect -8518 25222 -8462 25278
rect -8462 25222 -8458 25278
rect -8522 25218 -8458 25222
rect -8397 25278 -8333 25282
rect -8397 25222 -8393 25278
rect -8393 25222 -8337 25278
rect -8337 25222 -8333 25278
rect -8397 25218 -8333 25222
rect -6917 25268 -6853 25272
rect -6917 25212 -6913 25268
rect -6913 25212 -6857 25268
rect -6857 25212 -6853 25268
rect -6917 25208 -6853 25212
rect -6792 25268 -6728 25272
rect -6792 25212 -6788 25268
rect -6788 25212 -6732 25268
rect -6732 25212 -6728 25268
rect -6792 25208 -6728 25212
rect -6667 25268 -6603 25272
rect -6667 25212 -6663 25268
rect -6663 25212 -6607 25268
rect -6607 25212 -6603 25268
rect -6667 25208 -6603 25212
rect -472 24623 -408 24627
rect -472 24567 -468 24623
rect -468 24567 -412 24623
rect -412 24567 -408 24623
rect -472 24563 -408 24567
rect -472 24498 -408 24502
rect -472 24442 -468 24498
rect -468 24442 -412 24498
rect -412 24442 -408 24498
rect -472 24438 -408 24442
rect -472 24373 -408 24377
rect -472 24317 -468 24373
rect -468 24317 -412 24373
rect -412 24317 -408 24373
rect -472 24313 -408 24317
rect -492 23433 -428 23437
rect -492 23377 -488 23433
rect -488 23377 -432 23433
rect -432 23377 -428 23433
rect -492 23373 -428 23377
rect -492 23308 -428 23312
rect -492 23252 -488 23308
rect -488 23252 -432 23308
rect -432 23252 -428 23308
rect -492 23248 -428 23252
rect -492 23183 -428 23187
rect -492 23127 -488 23183
rect -488 23127 -432 23183
rect -432 23127 -428 23183
rect -492 23123 -428 23127
rect 963 23268 1027 23272
rect 963 23212 967 23268
rect 967 23212 1023 23268
rect 1023 23212 1027 23268
rect 963 23208 1027 23212
rect 1088 23268 1152 23272
rect 1088 23212 1092 23268
rect 1092 23212 1148 23268
rect 1148 23212 1152 23268
rect 1088 23208 1152 23212
rect 1213 23268 1277 23272
rect 1213 23212 1217 23268
rect 1217 23212 1273 23268
rect 1273 23212 1277 23268
rect 1213 23208 1277 23212
rect 1833 23278 1897 23282
rect 1833 23222 1837 23278
rect 1837 23222 1893 23278
rect 1893 23222 1897 23278
rect 1833 23218 1897 23222
rect 1958 23278 2022 23282
rect 1958 23222 1962 23278
rect 1962 23222 2018 23278
rect 2018 23222 2022 23278
rect 1958 23218 2022 23222
rect 2083 23278 2147 23282
rect 2083 23222 2087 23278
rect 2087 23222 2143 23278
rect 2143 23222 2147 23278
rect 2083 23218 2147 23222
rect 2733 23278 2797 23282
rect 2733 23222 2737 23278
rect 2737 23222 2793 23278
rect 2793 23222 2797 23278
rect 2733 23218 2797 23222
rect 2858 23278 2922 23282
rect 2858 23222 2862 23278
rect 2862 23222 2918 23278
rect 2918 23222 2922 23278
rect 2858 23218 2922 23222
rect 2983 23278 3047 23282
rect 2983 23222 2987 23278
rect 2987 23222 3043 23278
rect 3043 23222 3047 23278
rect 2983 23218 3047 23222
rect 3633 23278 3697 23282
rect 3633 23222 3637 23278
rect 3637 23222 3693 23278
rect 3693 23222 3697 23278
rect 3633 23218 3697 23222
rect 3758 23278 3822 23282
rect 3758 23222 3762 23278
rect 3762 23222 3818 23278
rect 3818 23222 3822 23278
rect 3758 23218 3822 23222
rect 3883 23278 3947 23282
rect 3883 23222 3887 23278
rect 3887 23222 3943 23278
rect 3943 23222 3947 23278
rect 3883 23218 3947 23222
rect 4523 23278 4587 23282
rect 4523 23222 4527 23278
rect 4527 23222 4583 23278
rect 4583 23222 4587 23278
rect 4523 23218 4587 23222
rect 4648 23278 4712 23282
rect 4648 23222 4652 23278
rect 4652 23222 4708 23278
rect 4708 23222 4712 23278
rect 4648 23218 4712 23222
rect 4773 23278 4837 23282
rect 4773 23222 4777 23278
rect 4777 23222 4833 23278
rect 4833 23222 4837 23278
rect 4773 23218 4837 23222
rect 5423 23278 5487 23282
rect 5423 23222 5427 23278
rect 5427 23222 5483 23278
rect 5483 23222 5487 23278
rect 5423 23218 5487 23222
rect 5548 23278 5612 23282
rect 5548 23222 5552 23278
rect 5552 23222 5608 23278
rect 5608 23222 5612 23278
rect 5548 23218 5612 23222
rect 5673 23278 5737 23282
rect 5673 23222 5677 23278
rect 5677 23222 5733 23278
rect 5733 23222 5737 23278
rect 5673 23218 5737 23222
rect 6333 23278 6397 23282
rect 6333 23222 6337 23278
rect 6337 23222 6393 23278
rect 6393 23222 6397 23278
rect 6333 23218 6397 23222
rect 6458 23278 6522 23282
rect 6458 23222 6462 23278
rect 6462 23222 6518 23278
rect 6518 23222 6522 23278
rect 6458 23218 6522 23222
rect 6583 23278 6647 23282
rect 6583 23222 6587 23278
rect 6587 23222 6643 23278
rect 6643 23222 6647 23278
rect 6583 23218 6647 23222
rect 6963 23278 7027 23282
rect 6963 23222 6967 23278
rect 6967 23222 7023 23278
rect 7023 23222 7027 23278
rect 6963 23218 7027 23222
rect 7088 23278 7152 23282
rect 7088 23222 7092 23278
rect 7092 23222 7148 23278
rect 7148 23222 7152 23278
rect 7088 23218 7152 23222
rect 7213 23278 7277 23282
rect 7213 23222 7217 23278
rect 7217 23222 7273 23278
rect 7273 23222 7277 23278
rect 7213 23218 7277 23222
rect 8153 23278 8217 23282
rect 8153 23222 8157 23278
rect 8157 23222 8213 23278
rect 8213 23222 8217 23278
rect 8153 23218 8217 23222
rect 8278 23278 8342 23282
rect 8278 23222 8282 23278
rect 8282 23222 8338 23278
rect 8338 23222 8342 23278
rect 8278 23218 8342 23222
rect 8403 23278 8467 23282
rect 8403 23222 8407 23278
rect 8407 23222 8463 23278
rect 8463 23222 8467 23278
rect 8403 23218 8467 23222
rect 9753 23278 9817 23282
rect 9753 23222 9757 23278
rect 9757 23222 9813 23278
rect 9813 23222 9817 23278
rect 9753 23218 9817 23222
rect 9878 23278 9942 23282
rect 9878 23222 9882 23278
rect 9882 23222 9938 23278
rect 9938 23222 9942 23278
rect 9878 23218 9942 23222
rect 10003 23278 10067 23282
rect 10003 23222 10007 23278
rect 10007 23222 10063 23278
rect 10063 23222 10067 23278
rect 10003 23218 10067 23222
rect 11323 23278 11387 23282
rect 11323 23222 11327 23278
rect 11327 23222 11383 23278
rect 11383 23222 11387 23278
rect 11323 23218 11387 23222
rect 11448 23278 11512 23282
rect 11448 23222 11452 23278
rect 11452 23222 11508 23278
rect 11508 23222 11512 23278
rect 11448 23218 11512 23222
rect 11573 23278 11637 23282
rect 11573 23222 11577 23278
rect 11577 23222 11633 23278
rect 11633 23222 11637 23278
rect 11573 23218 11637 23222
rect 13043 23278 13107 23282
rect 13043 23222 13047 23278
rect 13047 23222 13103 23278
rect 13103 23222 13107 23278
rect 13043 23218 13107 23222
rect 13168 23278 13232 23282
rect 13168 23222 13172 23278
rect 13172 23222 13228 23278
rect 13228 23222 13232 23278
rect 13168 23218 13232 23222
rect 13293 23278 13357 23282
rect 13293 23222 13297 23278
rect 13297 23222 13353 23278
rect 13353 23222 13357 23278
rect 13293 23218 13357 23222
rect 15853 23268 15917 23272
rect 15853 23212 15857 23268
rect 15857 23212 15913 23268
rect 15913 23212 15917 23268
rect 15853 23208 15917 23212
rect 15978 23268 16042 23272
rect 15978 23212 15982 23268
rect 15982 23212 16038 23268
rect 16038 23212 16042 23268
rect 15978 23208 16042 23212
rect 16103 23268 16167 23272
rect 16103 23212 16107 23268
rect 16107 23212 16163 23268
rect 16163 23212 16167 23268
rect 16103 23208 16167 23212
rect 19413 23268 19477 23272
rect 19413 23212 19417 23268
rect 19417 23212 19473 23268
rect 19473 23212 19477 23268
rect 19413 23208 19477 23212
rect 19538 23268 19602 23272
rect 19538 23212 19542 23268
rect 19542 23212 19598 23268
rect 19598 23212 19602 23268
rect 19538 23208 19602 23212
rect 19663 23268 19727 23272
rect 19663 23212 19667 23268
rect 19667 23212 19723 23268
rect 19723 23212 19727 23268
rect 19663 23208 19727 23212
rect 22693 23268 22757 23272
rect 22693 23212 22697 23268
rect 22697 23212 22753 23268
rect 22753 23212 22757 23268
rect 22693 23208 22757 23212
rect 22818 23268 22882 23272
rect 22818 23212 22822 23268
rect 22822 23212 22878 23268
rect 22878 23212 22882 23268
rect 22818 23208 22882 23212
rect 22943 23268 23007 23272
rect 22943 23212 22947 23268
rect 22947 23212 23003 23268
rect 23003 23212 23007 23268
rect 22943 23208 23007 23212
rect -10607 12718 -10543 12782
rect 23238 19523 23302 19527
rect 23238 19467 23242 19523
rect 23242 19467 23298 19523
rect 23298 19467 23302 19523
rect 23238 19463 23302 19467
rect 12608 19333 12672 19337
rect 12608 19277 12612 19333
rect 12612 19277 12668 19333
rect 12668 19277 12672 19333
rect 12608 19273 12672 19277
rect 12608 19208 12672 19212
rect 12608 19152 12612 19208
rect 12612 19152 12668 19208
rect 12668 19152 12672 19208
rect 12608 19148 12672 19152
rect 23238 19398 23302 19402
rect 23238 19342 23242 19398
rect 23242 19342 23298 19398
rect 23298 19342 23302 19398
rect 23238 19338 23302 19342
rect 23238 19273 23302 19277
rect 23238 19217 23242 19273
rect 23242 19217 23298 19273
rect 23298 19217 23302 19273
rect 23238 19213 23302 19217
rect 12608 19083 12672 19087
rect 12608 19027 12612 19083
rect 12612 19027 12668 19083
rect 12668 19027 12672 19083
rect 12608 19023 12672 19027
rect 12608 18603 12672 18607
rect 12608 18547 12612 18603
rect 12612 18547 12668 18603
rect 12668 18547 12672 18603
rect 12608 18543 12672 18547
rect 12608 18478 12672 18482
rect 12608 18422 12612 18478
rect 12612 18422 12668 18478
rect 12668 18422 12672 18478
rect 12608 18418 12672 18422
rect 11073 18358 11137 18362
rect 11073 18302 11077 18358
rect 11077 18302 11133 18358
rect 11133 18302 11137 18358
rect 11073 18298 11137 18302
rect 11198 18358 11262 18362
rect 11198 18302 11202 18358
rect 11202 18302 11258 18358
rect 11258 18302 11262 18358
rect 11198 18298 11262 18302
rect 12608 18353 12672 18357
rect 12608 18297 12612 18353
rect 12612 18297 12668 18353
rect 12668 18297 12672 18353
rect 12608 18293 12672 18297
rect 12513 18028 12577 18092
rect 12513 17198 12577 17262
rect 12513 15638 12577 15702
rect 12513 15448 12577 15512
rect 12703 17608 12767 17672
rect 14598 16168 14662 16172
rect 14598 16112 14602 16168
rect 14602 16112 14658 16168
rect 14658 16112 14662 16168
rect 14598 16108 14662 16112
rect 14598 16048 14662 16052
rect 14598 15992 14602 16048
rect 14602 15992 14658 16048
rect 14658 15992 14662 16048
rect 14598 15988 14662 15992
rect 23848 16068 23912 16132
rect 23968 16068 24032 16132
rect 29518 16112 29522 16132
rect 29522 16112 29578 16132
rect 29578 16112 29582 16132
rect 29518 16088 29582 16112
rect 29518 16068 29522 16088
rect 29522 16068 29578 16088
rect 29578 16068 29582 16088
rect 15098 15908 15162 15912
rect 15098 15852 15102 15908
rect 15102 15852 15158 15908
rect 15158 15852 15162 15908
rect 15098 15848 15162 15852
rect 15098 15788 15162 15792
rect 15098 15732 15102 15788
rect 15102 15732 15158 15788
rect 15158 15732 15162 15788
rect 15098 15728 15162 15732
rect 12583 15238 12647 15302
rect 12713 15238 12777 15302
rect 12583 15158 12647 15222
rect 12713 15158 12777 15222
rect -462 14988 -398 15052
rect -282 14988 -218 15052
rect -462 14808 -398 14872
rect -282 14808 -218 14872
rect -6982 12908 -6918 12912
rect -6982 12852 -6978 12908
rect -6978 12852 -6922 12908
rect -6922 12852 -6918 12908
rect -6982 12848 -6918 12852
rect -7352 12768 -7288 12772
rect -7352 12712 -7348 12768
rect -7348 12712 -7292 12768
rect -7292 12712 -7288 12768
rect -7352 12708 -7288 12712
rect -5402 12478 -5338 12542
rect -5282 12478 -5218 12542
rect -6582 11458 -6518 11462
rect -6582 11402 -6578 11458
rect -6578 11402 -6522 11458
rect -6522 11402 -6518 11458
rect -6582 11398 -6518 11402
rect -6462 11458 -6398 11462
rect -6462 11402 -6458 11458
rect -6458 11402 -6402 11458
rect -6402 11402 -6398 11458
rect -6462 11398 -6398 11402
rect -7312 11158 -7248 11222
rect -7192 11158 -7128 11222
rect -5822 10978 -5758 11042
rect -5702 10978 -5638 11042
rect -5222 12298 -5158 12362
rect -5102 12298 -5038 12362
rect -5222 10798 -5158 10862
rect -5042 12108 -4978 12172
rect -4922 12108 -4858 12172
rect -5162 10608 -5098 10672
rect -5042 10608 -4978 10672
rect 893 14988 957 14992
rect 893 14932 897 14988
rect 897 14932 953 14988
rect 953 14932 957 14988
rect 893 14928 957 14932
rect 1018 14988 1082 14992
rect 1018 14932 1022 14988
rect 1022 14932 1078 14988
rect 1078 14932 1082 14988
rect 1018 14928 1082 14932
rect 1143 14988 1207 14992
rect 1143 14932 1147 14988
rect 1147 14932 1203 14988
rect 1203 14932 1207 14988
rect 1143 14928 1207 14932
rect 893 14868 957 14872
rect 893 14812 897 14868
rect 897 14812 953 14868
rect 953 14812 957 14868
rect 893 14808 957 14812
rect 1018 14868 1082 14872
rect 1018 14812 1022 14868
rect 1022 14812 1078 14868
rect 1078 14812 1082 14868
rect 1018 14808 1082 14812
rect 1143 14868 1207 14872
rect 1143 14812 1147 14868
rect 1147 14812 1203 14868
rect 1203 14812 1207 14868
rect 1143 14808 1207 14812
rect 2613 14988 2677 14992
rect 2613 14932 2617 14988
rect 2617 14932 2673 14988
rect 2673 14932 2677 14988
rect 2613 14928 2677 14932
rect 2738 14988 2802 14992
rect 2738 14932 2742 14988
rect 2742 14932 2798 14988
rect 2798 14932 2802 14988
rect 2738 14928 2802 14932
rect 2863 14988 2927 14992
rect 2863 14932 2867 14988
rect 2867 14932 2923 14988
rect 2923 14932 2927 14988
rect 2863 14928 2927 14932
rect 2613 14868 2677 14872
rect 2613 14812 2617 14868
rect 2617 14812 2673 14868
rect 2673 14812 2677 14868
rect 2613 14808 2677 14812
rect 2738 14868 2802 14872
rect 2738 14812 2742 14868
rect 2742 14812 2798 14868
rect 2798 14812 2802 14868
rect 2738 14808 2802 14812
rect 2863 14868 2927 14872
rect 2863 14812 2867 14868
rect 2867 14812 2923 14868
rect 2923 14812 2927 14868
rect 2863 14808 2927 14812
rect 4053 14988 4117 14992
rect 4053 14932 4057 14988
rect 4057 14932 4113 14988
rect 4113 14932 4117 14988
rect 4053 14928 4117 14932
rect 4178 14988 4242 14992
rect 4178 14932 4182 14988
rect 4182 14932 4238 14988
rect 4238 14932 4242 14988
rect 4178 14928 4242 14932
rect 4303 14988 4367 14992
rect 4303 14932 4307 14988
rect 4307 14932 4363 14988
rect 4363 14932 4367 14988
rect 4303 14928 4367 14932
rect 4053 14868 4117 14872
rect 4053 14812 4057 14868
rect 4057 14812 4113 14868
rect 4113 14812 4117 14868
rect 4053 14808 4117 14812
rect 4178 14868 4242 14872
rect 4178 14812 4182 14868
rect 4182 14812 4238 14868
rect 4238 14812 4242 14868
rect 4178 14808 4242 14812
rect 4303 14868 4367 14872
rect 4303 14812 4307 14868
rect 4307 14812 4363 14868
rect 4363 14812 4367 14868
rect 4303 14808 4367 14812
rect 5513 14988 5577 14992
rect 5513 14932 5517 14988
rect 5517 14932 5573 14988
rect 5573 14932 5577 14988
rect 5513 14928 5577 14932
rect 5638 14988 5702 14992
rect 5638 14932 5642 14988
rect 5642 14932 5698 14988
rect 5698 14932 5702 14988
rect 5638 14928 5702 14932
rect 5763 14988 5827 14992
rect 5763 14932 5767 14988
rect 5767 14932 5823 14988
rect 5823 14932 5827 14988
rect 5763 14928 5827 14932
rect 5513 14868 5577 14872
rect 5513 14812 5517 14868
rect 5517 14812 5573 14868
rect 5573 14812 5577 14868
rect 5513 14808 5577 14812
rect 5638 14868 5702 14872
rect 5638 14812 5642 14868
rect 5642 14812 5698 14868
rect 5698 14812 5702 14868
rect 5638 14808 5702 14812
rect 5763 14868 5827 14872
rect 5763 14812 5767 14868
rect 5767 14812 5823 14868
rect 5823 14812 5827 14868
rect 5763 14808 5827 14812
rect 7353 14948 7417 14952
rect 7353 14892 7357 14948
rect 7357 14892 7413 14948
rect 7413 14892 7417 14948
rect 7353 14888 7417 14892
rect 7478 14948 7542 14952
rect 7478 14892 7482 14948
rect 7482 14892 7538 14948
rect 7538 14892 7542 14948
rect 7478 14888 7542 14892
rect 7603 14948 7667 14952
rect 7603 14892 7607 14948
rect 7607 14892 7663 14948
rect 7663 14892 7667 14948
rect 7603 14888 7667 14892
rect 8823 14958 8887 14962
rect 8823 14902 8827 14958
rect 8827 14902 8883 14958
rect 8883 14902 8887 14958
rect 8823 14898 8887 14902
rect 8948 14958 9012 14962
rect 8948 14902 8952 14958
rect 8952 14902 9008 14958
rect 9008 14902 9012 14958
rect 8948 14898 9012 14902
rect 9073 14958 9137 14962
rect 9073 14902 9077 14958
rect 9077 14902 9133 14958
rect 9133 14902 9137 14958
rect 9073 14898 9137 14902
rect 11683 14968 11747 14972
rect 11683 14912 11687 14968
rect 11687 14912 11743 14968
rect 11743 14912 11747 14968
rect 11683 14908 11747 14912
rect 11808 14968 11872 14972
rect 11808 14912 11812 14968
rect 11812 14912 11868 14968
rect 11868 14912 11872 14968
rect 11808 14908 11872 14912
rect 11933 14968 11997 14972
rect 11933 14912 11937 14968
rect 11937 14912 11993 14968
rect 11993 14912 11997 14968
rect 11933 14908 11997 14912
rect 12693 14968 12757 14972
rect 12693 14912 12697 14968
rect 12697 14912 12753 14968
rect 12753 14912 12757 14968
rect 12693 14908 12757 14912
rect 12818 14968 12882 14972
rect 12818 14912 12822 14968
rect 12822 14912 12878 14968
rect 12878 14912 12882 14968
rect 12818 14908 12882 14912
rect 12943 14968 13007 14972
rect 12943 14912 12947 14968
rect 12947 14912 13003 14968
rect 13003 14912 13007 14968
rect 12943 14908 13007 14912
rect 15263 14968 15327 14972
rect 15263 14912 15267 14968
rect 15267 14912 15323 14968
rect 15323 14912 15327 14968
rect 15263 14908 15327 14912
rect 15388 14968 15452 14972
rect 15388 14912 15392 14968
rect 15392 14912 15448 14968
rect 15448 14912 15452 14968
rect 15388 14908 15452 14912
rect 15513 14968 15577 14972
rect 15513 14912 15517 14968
rect 15517 14912 15573 14968
rect 15573 14912 15577 14968
rect 15513 14908 15577 14912
rect 15743 14968 15807 14972
rect 15743 14912 15747 14968
rect 15747 14912 15803 14968
rect 15803 14912 15807 14968
rect 15743 14908 15807 14912
rect 15868 14968 15932 14972
rect 15868 14912 15872 14968
rect 15872 14912 15928 14968
rect 15928 14912 15932 14968
rect 15868 14908 15932 14912
rect 15993 14968 16057 14972
rect 15993 14912 15997 14968
rect 15997 14912 16053 14968
rect 16053 14912 16057 14968
rect 15993 14908 16057 14912
rect 20523 14948 20587 14952
rect 20523 14892 20527 14948
rect 20527 14892 20583 14948
rect 20583 14892 20587 14948
rect 20523 14888 20587 14892
rect 20648 14948 20712 14952
rect 20648 14892 20652 14948
rect 20652 14892 20708 14948
rect 20708 14892 20712 14948
rect 20648 14888 20712 14892
rect 20773 14948 20837 14952
rect 20773 14892 20777 14948
rect 20777 14892 20833 14948
rect 20833 14892 20837 14948
rect 20773 14888 20837 14892
rect 20883 14948 20947 14952
rect 20883 14892 20887 14948
rect 20887 14892 20943 14948
rect 20943 14892 20947 14948
rect 20883 14888 20947 14892
rect 21008 14948 21072 14952
rect 21008 14892 21012 14948
rect 21012 14892 21068 14948
rect 21068 14892 21072 14948
rect 21008 14888 21072 14892
rect 21133 14948 21197 14952
rect 21133 14892 21137 14948
rect 21137 14892 21193 14948
rect 21193 14892 21197 14948
rect 21133 14888 21197 14892
rect 16088 14528 16152 14532
rect 16088 14472 16092 14528
rect 16092 14472 16148 14528
rect 16148 14472 16152 14528
rect 16088 14468 16152 14472
rect 20268 14528 20332 14532
rect 20268 14472 20272 14528
rect 20272 14472 20328 14528
rect 20328 14472 20332 14528
rect 20268 14468 20332 14472
rect 23968 14318 24032 14382
rect 22308 14198 22372 14202
rect 22308 14142 22312 14198
rect 22312 14142 22368 14198
rect 22368 14142 22372 14198
rect 22308 14138 22372 14142
rect 23968 14198 24032 14262
rect 24168 15808 24232 15872
rect 24288 15808 24352 15872
rect 29338 15852 29342 15872
rect 29342 15852 29398 15872
rect 29398 15852 29402 15872
rect 29338 15828 29402 15852
rect 29338 15808 29342 15828
rect 29342 15808 29398 15828
rect 29398 15808 29402 15828
rect 26763 15478 26827 15542
rect 26863 15478 26927 15542
rect 26523 15198 26587 15262
rect 26623 15198 26687 15262
rect 24168 14318 24232 14382
rect 24168 14198 24232 14262
rect 26828 14313 26892 14377
rect 258 13778 322 13842
rect 378 13778 442 13842
rect 138 12478 202 12542
rect 258 12478 322 12542
rect 438 13598 502 13662
rect 558 13598 622 13662
rect 318 12298 382 12362
rect 438 12298 502 12362
rect 618 13408 682 13472
rect 738 13408 802 13472
rect 498 12108 562 12172
rect 618 12108 682 12172
rect -442 11398 -378 11462
rect -312 11398 -248 11462
rect -5522 10428 -5458 10492
rect -5402 10428 -5338 10492
rect -5707 8928 -5643 8992
rect -5577 8928 -5513 8992
rect 263 8928 327 8992
rect 393 8928 457 8992
rect -462 7508 -398 7572
rect -282 7508 -218 7572
rect -462 7328 -398 7392
rect -282 7328 -218 7392
rect -6567 923 -6503 987
rect -6447 923 -6383 987
rect -6077 913 -6013 977
rect -5947 913 -5883 977
rect 953 7478 1017 7482
rect 953 7422 957 7478
rect 957 7422 1013 7478
rect 1013 7422 1017 7478
rect 953 7418 1017 7422
rect 1078 7478 1142 7482
rect 1078 7422 1082 7478
rect 1082 7422 1138 7478
rect 1138 7422 1142 7478
rect 1078 7418 1142 7422
rect 1563 7478 1627 7482
rect 1563 7422 1567 7478
rect 1567 7422 1623 7478
rect 1623 7422 1627 7478
rect 1563 7418 1627 7422
rect 1688 7478 1752 7482
rect 1688 7422 1692 7478
rect 1692 7422 1748 7478
rect 1748 7422 1752 7478
rect 1688 7418 1752 7422
rect 2713 7478 2777 7482
rect 2713 7422 2717 7478
rect 2717 7422 2773 7478
rect 2773 7422 2777 7478
rect 2713 7418 2777 7422
rect 2838 7478 2902 7482
rect 2838 7422 2842 7478
rect 2842 7422 2898 7478
rect 2898 7422 2902 7478
rect 2838 7418 2902 7422
rect 3883 7478 3947 7482
rect 3883 7422 3887 7478
rect 3887 7422 3943 7478
rect 3943 7422 3947 7478
rect 3883 7418 3947 7422
rect 4008 7478 4072 7482
rect 4008 7422 4012 7478
rect 4012 7422 4068 7478
rect 4068 7422 4072 7478
rect 4008 7418 4072 7422
rect 5043 7478 5107 7482
rect 5043 7422 5047 7478
rect 5047 7422 5103 7478
rect 5103 7422 5107 7478
rect 5043 7418 5107 7422
rect 5168 7478 5232 7482
rect 5168 7422 5172 7478
rect 5172 7422 5228 7478
rect 5228 7422 5232 7478
rect 5168 7418 5232 7422
rect 6213 7478 6277 7482
rect 6213 7422 6217 7478
rect 6217 7422 6273 7478
rect 6273 7422 6277 7478
rect 6213 7418 6277 7422
rect 6338 7478 6402 7482
rect 6338 7422 6342 7478
rect 6342 7422 6398 7478
rect 6398 7422 6402 7478
rect 6338 7418 6402 7422
rect 7373 7478 7437 7482
rect 7373 7422 7377 7478
rect 7377 7422 7433 7478
rect 7433 7422 7437 7478
rect 7373 7418 7437 7422
rect 7498 7478 7562 7482
rect 7498 7422 7502 7478
rect 7502 7422 7558 7478
rect 7558 7422 7562 7478
rect 7498 7418 7562 7422
rect 373 6748 437 6812
rect 483 6748 547 6812
rect 22308 3893 22372 3957
rect -462 408 -398 472
rect -282 408 -218 472
rect 1393 408 1457 412
rect 1393 352 1397 408
rect 1397 352 1453 408
rect 1453 352 1457 408
rect 1393 348 1457 352
rect 1518 408 1582 412
rect 1518 352 1522 408
rect 1522 352 1578 408
rect 1578 352 1582 408
rect 1518 348 1582 352
rect 1643 408 1707 412
rect 1643 352 1647 408
rect 1647 352 1703 408
rect 1703 352 1707 408
rect 1643 348 1707 352
rect 3123 408 3187 412
rect 3123 352 3127 408
rect 3127 352 3183 408
rect 3183 352 3187 408
rect 3123 348 3187 352
rect 3248 408 3312 412
rect 3248 352 3252 408
rect 3252 352 3308 408
rect 3308 352 3312 408
rect 3248 348 3312 352
rect 3373 408 3437 412
rect 3373 352 3377 408
rect 3377 352 3433 408
rect 3433 352 3437 408
rect 3373 348 3437 352
rect 5183 408 5247 412
rect 5183 352 5187 408
rect 5187 352 5243 408
rect 5243 352 5247 408
rect 5183 348 5247 352
rect 5308 408 5372 412
rect 5308 352 5312 408
rect 5312 352 5368 408
rect 5368 352 5372 408
rect 5308 348 5372 352
rect 5433 408 5497 412
rect 5433 352 5437 408
rect 5437 352 5493 408
rect 5493 352 5497 408
rect 5433 348 5497 352
rect 8823 398 8887 402
rect 8823 342 8827 398
rect 8827 342 8883 398
rect 8883 342 8887 398
rect 8823 338 8887 342
rect 8948 398 9012 402
rect 8948 342 8952 398
rect 8952 342 9008 398
rect 9008 342 9012 398
rect 8948 338 9012 342
rect 9073 398 9137 402
rect 9073 342 9077 398
rect 9077 342 9133 398
rect 9133 342 9137 398
rect 9073 338 9137 342
rect 10943 398 11007 402
rect 10943 342 10947 398
rect 10947 342 11003 398
rect 11003 342 11007 398
rect 10943 338 11007 342
rect 11068 398 11132 402
rect 11068 342 11072 398
rect 11072 342 11128 398
rect 11128 342 11132 398
rect 11068 338 11132 342
rect 11193 398 11257 402
rect 11193 342 11197 398
rect 11197 342 11253 398
rect 11253 342 11257 398
rect 11193 338 11257 342
rect 14673 398 14737 402
rect 14673 342 14677 398
rect 14677 342 14733 398
rect 14733 342 14737 398
rect 14673 338 14737 342
rect 14798 398 14862 402
rect 14798 342 14802 398
rect 14802 342 14858 398
rect 14858 342 14862 398
rect 14798 338 14862 342
rect 14923 398 14987 402
rect 14923 342 14927 398
rect 14927 342 14983 398
rect 14983 342 14987 398
rect 14923 338 14987 342
rect 17033 398 17097 402
rect 17033 342 17037 398
rect 17037 342 17093 398
rect 17093 342 17097 398
rect 17033 338 17097 342
rect 17158 398 17222 402
rect 17158 342 17162 398
rect 17162 342 17218 398
rect 17218 342 17222 398
rect 17158 338 17222 342
rect 17283 398 17347 402
rect 17283 342 17287 398
rect 17287 342 17343 398
rect 17343 342 17347 398
rect 17283 338 17347 342
rect 19043 398 19107 402
rect 19043 342 19047 398
rect 19047 342 19103 398
rect 19103 342 19107 398
rect 19043 338 19107 342
rect 19168 398 19232 402
rect 19168 342 19172 398
rect 19172 342 19228 398
rect 19228 342 19232 398
rect 19168 338 19232 342
rect 19293 398 19357 402
rect 19293 342 19297 398
rect 19297 342 19353 398
rect 19353 342 19357 398
rect 19293 338 19357 342
rect 21003 398 21067 402
rect 21003 342 21007 398
rect 21007 342 21063 398
rect 21063 342 21067 398
rect 21003 338 21067 342
rect 21128 398 21192 402
rect 21128 342 21132 398
rect 21132 342 21188 398
rect 21188 342 21192 398
rect 21128 338 21192 342
rect 21253 398 21317 402
rect 21253 342 21257 398
rect 21257 342 21313 398
rect 21313 342 21317 398
rect 21253 338 21317 342
rect -462 228 -398 292
rect -282 228 -218 292
<< metal4 >>
rect -10950 25282 -220 25380
rect -10950 25272 -8647 25282
rect -10950 25208 -10417 25272
rect -10353 25208 -10292 25272
rect -10228 25208 -10167 25272
rect -10103 25218 -8647 25272
rect -8583 25218 -8522 25282
rect -8458 25218 -8397 25282
rect -8333 25272 -220 25282
rect -8333 25218 -6917 25272
rect -10103 25208 -6917 25218
rect -6853 25208 -6792 25272
rect -6728 25208 -6667 25272
rect -6603 25208 -220 25272
rect -10950 25080 -220 25208
rect -520 24627 -220 25080
rect -520 24563 -472 24627
rect -408 24563 -220 24627
rect -520 24502 -220 24563
rect -520 24438 -472 24502
rect -408 24438 -220 24502
rect -520 24377 -220 24438
rect -520 24313 -472 24377
rect -408 24313 -220 24377
rect -520 23437 -220 24313
rect -520 23373 -492 23437
rect -428 23400 -220 23437
rect -428 23373 23510 23400
rect -520 23312 23510 23373
rect -520 23248 -492 23312
rect -428 23282 23510 23312
rect -428 23272 1833 23282
rect -428 23248 963 23272
rect -520 23208 963 23248
rect 1027 23208 1088 23272
rect 1152 23208 1213 23272
rect 1277 23218 1833 23272
rect 1897 23218 1958 23282
rect 2022 23218 2083 23282
rect 2147 23218 2733 23282
rect 2797 23218 2858 23282
rect 2922 23218 2983 23282
rect 3047 23218 3633 23282
rect 3697 23218 3758 23282
rect 3822 23218 3883 23282
rect 3947 23218 4523 23282
rect 4587 23218 4648 23282
rect 4712 23218 4773 23282
rect 4837 23218 5423 23282
rect 5487 23218 5548 23282
rect 5612 23218 5673 23282
rect 5737 23218 6333 23282
rect 6397 23218 6458 23282
rect 6522 23218 6583 23282
rect 6647 23218 6963 23282
rect 7027 23218 7088 23282
rect 7152 23218 7213 23282
rect 7277 23218 8153 23282
rect 8217 23218 8278 23282
rect 8342 23218 8403 23282
rect 8467 23218 9753 23282
rect 9817 23218 9878 23282
rect 9942 23218 10003 23282
rect 10067 23218 11323 23282
rect 11387 23218 11448 23282
rect 11512 23218 11573 23282
rect 11637 23218 13043 23282
rect 13107 23218 13168 23282
rect 13232 23218 13293 23282
rect 13357 23272 23510 23282
rect 13357 23218 15853 23272
rect 1277 23208 15853 23218
rect 15917 23208 15978 23272
rect 16042 23208 16103 23272
rect 16167 23208 19413 23272
rect 19477 23208 19538 23272
rect 19602 23208 19663 23272
rect 19727 23208 22693 23272
rect 22757 23208 22818 23272
rect 22882 23208 22943 23272
rect 23007 23208 23510 23272
rect -520 23187 23510 23208
rect -520 23123 -492 23187
rect -428 23123 23510 23187
rect -520 23100 23510 23123
rect 12490 19337 12790 23100
rect 12490 19273 12608 19337
rect 12672 19273 12790 19337
rect 12490 19212 12790 19273
rect 12490 19148 12608 19212
rect 12672 19148 12790 19212
rect 23210 19527 23510 23100
rect 23210 19463 23238 19527
rect 23302 19463 23510 19527
rect 23210 19402 23510 19463
rect 23210 19338 23238 19402
rect 23302 19338 23510 19402
rect 23210 19277 23510 19338
rect 23210 19213 23238 19277
rect 23302 19213 23510 19277
rect 23210 19190 23510 19213
rect 12490 19087 12790 19148
rect 12490 19023 12608 19087
rect 12672 19023 12790 19087
rect 12490 18607 12790 19023
rect 12490 18543 12608 18607
rect 12672 18543 12790 18607
rect 12490 18490 12790 18543
rect 11000 18482 12790 18490
rect 11000 18418 12608 18482
rect 12672 18418 12790 18482
rect 11000 18362 12790 18418
rect 11000 18298 11073 18362
rect 11137 18298 11198 18362
rect 11262 18357 12790 18362
rect 11262 18298 12608 18357
rect 11000 18293 12608 18298
rect 12672 18293 12790 18357
rect 11000 18190 12790 18293
rect 12480 18092 12670 18110
rect 12480 18028 12513 18092
rect 12577 18030 12670 18092
rect 12577 18028 12610 18030
rect 12480 18010 12610 18028
rect 12670 17672 12800 17690
rect 12670 17608 12703 17672
rect 12767 17608 12800 17672
rect 12670 17590 12800 17608
rect 12480 17270 12610 17280
rect 12480 17262 12800 17270
rect 12480 17198 12513 17262
rect 12577 17198 12800 17262
rect 12480 17190 12800 17198
rect 12480 17180 12610 17190
rect 29930 16190 30230 16310
rect 14580 16172 30230 16190
rect 14580 16108 14598 16172
rect 14662 16132 30230 16172
rect 14662 16108 23848 16132
rect 14580 16068 23848 16108
rect 23912 16068 23968 16132
rect 24032 16068 29518 16132
rect 29582 16068 30230 16132
rect 14580 16052 30230 16068
rect 14580 15988 14598 16052
rect 14662 16010 30230 16052
rect 14662 15988 14680 16010
rect 14580 15970 14680 15988
rect 15080 15912 30050 15930
rect 15080 15848 15098 15912
rect 15162 15872 30050 15912
rect 15162 15848 24168 15872
rect 15080 15808 24168 15848
rect 24232 15808 24288 15872
rect 24352 15808 29338 15872
rect 29402 15808 30050 15872
rect 15080 15792 30050 15808
rect 12480 15730 12600 15731
rect 12480 15702 12610 15730
rect 15080 15728 15098 15792
rect 15162 15750 30050 15792
rect 15162 15728 15180 15750
rect 15080 15710 15180 15728
rect 12480 15638 12513 15702
rect 12577 15638 12610 15702
rect 12480 15600 12610 15638
rect 30310 15630 30610 15930
rect 12480 15542 26940 15600
rect 12480 15512 26763 15542
rect 12480 15448 12513 15512
rect 12577 15478 26763 15512
rect 26827 15478 26863 15542
rect 26927 15478 26940 15542
rect 12577 15448 26940 15478
rect 12480 15420 26940 15448
rect 12510 15302 26701 15320
rect 12510 15238 12583 15302
rect 12647 15238 12713 15302
rect 12777 15262 26701 15302
rect 12777 15238 26523 15262
rect 12510 15222 26523 15238
rect 12510 15158 12583 15222
rect 12647 15158 12713 15222
rect 12777 15198 26523 15222
rect 26587 15198 26623 15262
rect 26687 15198 26701 15262
rect 12777 15158 26701 15198
rect 12510 15140 26701 15158
rect -490 15052 23760 15080
rect -490 14988 -462 15052
rect -398 14988 -282 15052
rect -218 14992 23760 15052
rect -218 14988 893 14992
rect -490 14928 893 14988
rect 957 14928 1018 14992
rect 1082 14928 1143 14992
rect 1207 14928 2613 14992
rect 2677 14928 2738 14992
rect 2802 14928 2863 14992
rect 2927 14928 4053 14992
rect 4117 14928 4178 14992
rect 4242 14928 4303 14992
rect 4367 14928 5513 14992
rect 5577 14928 5638 14992
rect 5702 14928 5763 14992
rect 5827 14972 23760 14992
rect 5827 14962 11683 14972
rect 5827 14952 8823 14962
rect 5827 14928 7353 14952
rect -490 14888 7353 14928
rect 7417 14888 7478 14952
rect 7542 14888 7603 14952
rect 7667 14898 8823 14952
rect 8887 14898 8948 14962
rect 9012 14898 9073 14962
rect 9137 14908 11683 14962
rect 11747 14908 11808 14972
rect 11872 14908 11933 14972
rect 11997 14908 12693 14972
rect 12757 14908 12818 14972
rect 12882 14908 12943 14972
rect 13007 14908 15263 14972
rect 15327 14908 15388 14972
rect 15452 14908 15513 14972
rect 15577 14908 15743 14972
rect 15807 14908 15868 14972
rect 15932 14908 15993 14972
rect 16057 14952 23760 14972
rect 16057 14908 20523 14952
rect 9137 14898 20523 14908
rect 7667 14888 20523 14898
rect 20587 14888 20648 14952
rect 20712 14888 20773 14952
rect 20837 14888 20883 14952
rect 20947 14888 21008 14952
rect 21072 14888 21133 14952
rect 21197 14888 23760 14952
rect -490 14872 23760 14888
rect -490 14808 -462 14872
rect -398 14808 -282 14872
rect -218 14808 893 14872
rect 957 14808 1018 14872
rect 1082 14808 1143 14872
rect 1207 14808 2613 14872
rect 2677 14808 2738 14872
rect 2802 14808 2863 14872
rect 2927 14808 4053 14872
rect 4117 14808 4178 14872
rect 4242 14808 4303 14872
rect 4367 14808 5513 14872
rect 5577 14808 5638 14872
rect 5702 14808 5763 14872
rect 5827 14808 23760 14872
rect -490 14780 23760 14808
rect 15500 14532 20350 14550
rect 15500 14470 16088 14532
rect 15500 14110 15580 14470
rect 16070 14468 16088 14470
rect 16152 14470 20268 14532
rect 16152 14468 16170 14470
rect 16070 14450 16170 14468
rect 20250 14468 20268 14470
rect 20332 14468 20350 14532
rect 20250 14450 20350 14468
rect 22280 14202 22400 14220
rect 22280 14138 22308 14202
rect 22372 14138 22400 14202
rect 230 13842 470 13870
rect 230 13778 258 13842
rect 322 13778 378 13842
rect 442 13778 470 13842
rect 230 13750 470 13778
rect 410 13662 650 13690
rect 410 13598 438 13662
rect 502 13598 558 13662
rect 622 13598 650 13662
rect 410 13570 650 13598
rect 590 13472 830 13500
rect 590 13408 618 13472
rect 682 13408 738 13472
rect 802 13408 830 13472
rect 590 13380 830 13408
rect -7450 12912 -6900 12930
rect -7450 12850 -6982 12912
rect -7000 12848 -6982 12850
rect -6918 12848 -6900 12912
rect -7000 12830 -6900 12848
rect -10620 12790 -10530 12800
rect -10620 12782 -7270 12790
rect -10620 12718 -10607 12782
rect -10543 12772 -7270 12782
rect -10543 12718 -7352 12772
rect -10620 12710 -7352 12718
rect -10620 12700 -10530 12710
rect -7370 12708 -7352 12710
rect -7288 12708 -7270 12772
rect -7370 12690 -7270 12708
rect -5430 12542 350 12570
rect -5430 12478 -5402 12542
rect -5338 12478 -5282 12542
rect -5218 12478 138 12542
rect 202 12478 258 12542
rect 322 12478 350 12542
rect -5430 12450 350 12478
rect -5250 12362 530 12390
rect -5250 12298 -5222 12362
rect -5158 12298 -5102 12362
rect -5038 12298 318 12362
rect 382 12298 438 12362
rect 502 12298 530 12362
rect -5250 12270 530 12298
rect -5070 12172 710 12200
rect -5070 12108 -5042 12172
rect -4978 12108 -4922 12172
rect -4858 12108 498 12172
rect 562 12108 618 12172
rect 682 12108 710 12172
rect -5070 12080 710 12108
rect -6600 11462 -190 11480
rect -6600 11398 -6582 11462
rect -6518 11398 -6462 11462
rect -6398 11398 -442 11462
rect -378 11398 -312 11462
rect -248 11398 -190 11462
rect -6600 11380 -190 11398
rect -10830 11250 -10530 11340
rect -10830 11222 -7110 11250
rect -10830 11158 -7312 11222
rect -7248 11158 -7192 11222
rect -7128 11158 -7110 11222
rect -10830 11130 -7110 11158
rect -10830 11040 -10530 11130
rect -9700 11042 -5610 11070
rect -9700 10978 -5822 11042
rect -5758 10978 -5702 11042
rect -5638 10978 -5610 11042
rect -9700 10950 -5610 10978
rect -9090 10862 -5130 10890
rect -9090 10798 -5222 10862
rect -5158 10798 -5130 10862
rect -9090 10770 -5130 10798
rect -1930 10810 -640 11000
rect -1930 10700 280 10810
rect -8500 10672 -4950 10700
rect -8500 10608 -5162 10672
rect -5098 10608 -5042 10672
rect -4978 10608 -4950 10672
rect -8500 10580 -4950 10608
rect -7920 10492 -5310 10520
rect -7920 10428 -5522 10492
rect -5458 10428 -5402 10492
rect -5338 10428 -5310 10492
rect -7920 10400 -5310 10428
rect -1930 10040 -1630 10700
rect -10840 9740 -1630 10040
rect -1350 10400 280 10510
rect -1350 10210 -640 10400
rect -1350 9500 -1050 10210
rect -10820 9200 -1050 9500
rect -5730 8992 480 9020
rect -5730 8928 -5707 8992
rect -5643 8928 -5577 8992
rect -5513 8928 263 8992
rect 327 8928 393 8992
rect 457 8928 480 8992
rect -5730 8900 480 8928
rect -490 7572 7620 7600
rect -490 7508 -462 7572
rect -398 7508 -282 7572
rect -218 7508 7620 7572
rect -490 7482 7620 7508
rect -490 7418 953 7482
rect 1017 7418 1078 7482
rect 1142 7418 1563 7482
rect 1627 7418 1688 7482
rect 1752 7418 2713 7482
rect 2777 7418 2838 7482
rect 2902 7418 3883 7482
rect 3947 7418 4008 7482
rect 4072 7418 5043 7482
rect 5107 7418 5168 7482
rect 5232 7418 6213 7482
rect 6277 7418 6338 7482
rect 6402 7418 7373 7482
rect 7437 7418 7498 7482
rect 7562 7418 7620 7482
rect -490 7392 7620 7418
rect -490 7328 -462 7392
rect -398 7328 -282 7392
rect -218 7328 7620 7392
rect -490 7300 7620 7328
rect 360 6812 560 6830
rect 360 6748 373 6812
rect 437 6748 483 6812
rect 547 6748 560 6812
rect 360 6730 560 6748
rect 22280 3957 22400 14138
rect 22630 13830 22730 14780
rect 23950 14382 24050 14400
rect 23950 14318 23968 14382
rect 24032 14318 24050 14382
rect 23950 14262 24050 14318
rect 23950 14198 23968 14262
rect 24032 14198 24050 14262
rect 23950 14180 24050 14198
rect 24150 14382 24250 14400
rect 24150 14318 24168 14382
rect 24232 14318 24250 14382
rect 24150 14262 24250 14318
rect 26810 14377 26910 14390
rect 26810 14313 26828 14377
rect 26892 14313 26910 14377
rect 26810 14300 26910 14313
rect 24150 14198 24168 14262
rect 24232 14198 24250 14262
rect 24150 14180 24250 14198
rect 22280 3893 22308 3957
rect 22372 3893 22400 3957
rect 22280 3870 22400 3893
rect -6570 987 -6500 1020
rect -6570 923 -6567 987
rect -6503 923 -6500 987
rect -6570 890 -6500 923
rect -6450 987 -6380 1020
rect -6450 923 -6447 987
rect -6383 923 -6380 987
rect -6450 890 -6380 923
rect -6110 977 -5860 1040
rect -6110 913 -6077 977
rect -6013 913 -5947 977
rect -5883 913 -5860 977
rect -6110 870 -5860 913
rect -11080 472 22730 490
rect -11080 408 -462 472
rect -398 408 -282 472
rect -218 412 22730 472
rect -218 408 1393 412
rect -11080 348 1393 408
rect 1457 348 1518 412
rect 1582 348 1643 412
rect 1707 348 3123 412
rect 3187 348 3248 412
rect 3312 348 3373 412
rect 3437 348 5183 412
rect 5247 348 5308 412
rect 5372 348 5433 412
rect 5497 402 22730 412
rect 5497 348 8823 402
rect -11080 338 8823 348
rect 8887 338 8948 402
rect 9012 338 9073 402
rect 9137 338 10943 402
rect 11007 338 11068 402
rect 11132 338 11193 402
rect 11257 338 14673 402
rect 14737 338 14798 402
rect 14862 338 14923 402
rect 14987 338 17033 402
rect 17097 338 17158 402
rect 17222 338 17283 402
rect 17347 338 19043 402
rect 19107 338 19168 402
rect 19232 338 19293 402
rect 19357 338 21003 402
rect 21067 338 21128 402
rect 21192 338 21253 402
rect 21317 338 22730 402
rect -11080 292 22730 338
rect -11080 228 -462 292
rect -398 228 -282 292
rect -218 228 22730 292
rect -11080 190 22730 228
rect 22190 -40 22490 130
rect -11080 -340 22490 -40
use bias_dummy  bias_dummy_0
timestamp 1757161594
transform 0 1 -1320 1 0 11100
box 1670 -8950 13960 750
use block01  block01_0
timestamp 1757161594
transform 1 0 14270 0 1 18790
box -1800 -2510 3461 80
use block03  block03_0
timestamp 1757161594
transform 0 -1 20200 -1 0 13850
box -790 -436 1246 4596
use block04  block04_0
timestamp 1757161594
transform 0 -1 20570 1 0 16850
box -570 -2970 2080 2840
use block02  block0102_0
timestamp 1757161594
transform 1 0 12780 0 1 17830
box -1196 -5226 2816 -2890
use cap  cap_1
timestamp 1757161594
transform 0 -1 31842 1 0 -1050
box 900 980 15510 9252
use cs_p_5  cs_p_5_0
timestamp 1757161594
transform 0 1 13293 1 0 19020
box -240 -413 4063 9820
use Diff_opamp_ly  Diff_opamp_ly_0
timestamp 1757161594
transform 1 0 -60 0 1 1230
box -60 -1230 22531 21951
use nmos_08  nmos_08_0
timestamp 1757161594
transform 0 -1 21986 1 0 12700
box 0 -26 1634 1212
use res  res_0
timestamp 1757161594
transform -1 0 29753 0 -1 25390
box -163 -193 6143 9070
use switchblock01  switchblock_0
timestamp 1757161594
transform 1 0 -10440 0 1 22920
box -628 -2220 4000 1868
use switchblock  switchblock_1
timestamp 1757161594
transform 0 -1 -9790 -1 0 11940
box -12993 -4583 1540 1123
<< end >>
