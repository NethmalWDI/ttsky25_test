magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -386 -669 386 669
<< nmoslvt >>
rect -200 -531 200 469
<< ndiff >>
rect -258 428 -200 469
rect -258 394 -246 428
rect -212 394 -200 428
rect -258 360 -200 394
rect -258 326 -246 360
rect -212 326 -200 360
rect -258 292 -200 326
rect -258 258 -246 292
rect -212 258 -200 292
rect -258 224 -200 258
rect -258 190 -246 224
rect -212 190 -200 224
rect -258 156 -200 190
rect -258 122 -246 156
rect -212 122 -200 156
rect -258 88 -200 122
rect -258 54 -246 88
rect -212 54 -200 88
rect -258 20 -200 54
rect -258 -14 -246 20
rect -212 -14 -200 20
rect -258 -48 -200 -14
rect -258 -82 -246 -48
rect -212 -82 -200 -48
rect -258 -116 -200 -82
rect -258 -150 -246 -116
rect -212 -150 -200 -116
rect -258 -184 -200 -150
rect -258 -218 -246 -184
rect -212 -218 -200 -184
rect -258 -252 -200 -218
rect -258 -286 -246 -252
rect -212 -286 -200 -252
rect -258 -320 -200 -286
rect -258 -354 -246 -320
rect -212 -354 -200 -320
rect -258 -388 -200 -354
rect -258 -422 -246 -388
rect -212 -422 -200 -388
rect -258 -456 -200 -422
rect -258 -490 -246 -456
rect -212 -490 -200 -456
rect -258 -531 -200 -490
rect 200 428 258 469
rect 200 394 212 428
rect 246 394 258 428
rect 200 360 258 394
rect 200 326 212 360
rect 246 326 258 360
rect 200 292 258 326
rect 200 258 212 292
rect 246 258 258 292
rect 200 224 258 258
rect 200 190 212 224
rect 246 190 258 224
rect 200 156 258 190
rect 200 122 212 156
rect 246 122 258 156
rect 200 88 258 122
rect 200 54 212 88
rect 246 54 258 88
rect 200 20 258 54
rect 200 -14 212 20
rect 246 -14 258 20
rect 200 -48 258 -14
rect 200 -82 212 -48
rect 246 -82 258 -48
rect 200 -116 258 -82
rect 200 -150 212 -116
rect 246 -150 258 -116
rect 200 -184 258 -150
rect 200 -218 212 -184
rect 246 -218 258 -184
rect 200 -252 258 -218
rect 200 -286 212 -252
rect 246 -286 258 -252
rect 200 -320 258 -286
rect 200 -354 212 -320
rect 246 -354 258 -320
rect 200 -388 258 -354
rect 200 -422 212 -388
rect 246 -422 258 -388
rect 200 -456 258 -422
rect 200 -490 212 -456
rect 246 -490 258 -456
rect 200 -531 258 -490
<< ndiffc >>
rect -246 394 -212 428
rect -246 326 -212 360
rect -246 258 -212 292
rect -246 190 -212 224
rect -246 122 -212 156
rect -246 54 -212 88
rect -246 -14 -212 20
rect -246 -82 -212 -48
rect -246 -150 -212 -116
rect -246 -218 -212 -184
rect -246 -286 -212 -252
rect -246 -354 -212 -320
rect -246 -422 -212 -388
rect -246 -490 -212 -456
rect 212 394 246 428
rect 212 326 246 360
rect 212 258 246 292
rect 212 190 246 224
rect 212 122 246 156
rect 212 54 246 88
rect 212 -14 246 20
rect 212 -82 246 -48
rect 212 -150 246 -116
rect 212 -218 246 -184
rect 212 -286 246 -252
rect 212 -354 246 -320
rect 212 -422 246 -388
rect 212 -490 246 -456
<< psubdiff >>
rect -360 609 360 643
rect -360 -609 -326 609
rect 326 -609 360 609
rect -360 -643 360 -609
<< poly >>
rect -200 541 200 557
rect -200 507 -153 541
rect -119 507 -85 541
rect -51 507 -17 541
rect 17 507 51 541
rect 85 507 119 541
rect 153 507 200 541
rect -200 469 200 507
rect -200 -557 200 -531
<< polycont >>
rect -153 507 -119 541
rect -85 507 -51 541
rect -17 507 17 541
rect 51 507 85 541
rect 119 507 153 541
<< locali >>
rect -360 609 360 643
rect -360 -609 -326 609
rect -200 507 -161 541
rect -119 507 -89 541
rect -51 507 -17 541
rect 17 507 51 541
rect 89 507 119 541
rect 161 507 200 541
rect -246 454 -212 473
rect -246 382 -212 394
rect -246 310 -212 326
rect -246 238 -212 258
rect -246 166 -212 190
rect -246 94 -212 122
rect -246 22 -212 54
rect -246 -48 -212 -14
rect -246 -116 -212 -84
rect -246 -184 -212 -156
rect -246 -252 -212 -228
rect -246 -320 -212 -300
rect -246 -388 -212 -372
rect -246 -456 -212 -444
rect -246 -535 -212 -516
rect 212 454 246 473
rect 212 382 246 394
rect 212 310 246 326
rect 212 238 246 258
rect 212 166 246 190
rect 212 94 246 122
rect 212 22 246 54
rect 212 -48 246 -14
rect 212 -116 246 -84
rect 212 -184 246 -156
rect 212 -252 246 -228
rect 212 -320 246 -300
rect 212 -388 246 -372
rect 212 -456 246 -444
rect 212 -535 246 -516
rect 326 -609 360 609
rect -360 -643 360 -609
<< viali >>
rect -161 507 -153 541
rect -153 507 -127 541
rect -89 507 -85 541
rect -85 507 -55 541
rect -17 507 17 541
rect 55 507 85 541
rect 85 507 89 541
rect 127 507 153 541
rect 153 507 161 541
rect -246 428 -212 454
rect -246 420 -212 428
rect -246 360 -212 382
rect -246 348 -212 360
rect -246 292 -212 310
rect -246 276 -212 292
rect -246 224 -212 238
rect -246 204 -212 224
rect -246 156 -212 166
rect -246 132 -212 156
rect -246 88 -212 94
rect -246 60 -212 88
rect -246 20 -212 22
rect -246 -12 -212 20
rect -246 -82 -212 -50
rect -246 -84 -212 -82
rect -246 -150 -212 -122
rect -246 -156 -212 -150
rect -246 -218 -212 -194
rect -246 -228 -212 -218
rect -246 -286 -212 -266
rect -246 -300 -212 -286
rect -246 -354 -212 -338
rect -246 -372 -212 -354
rect -246 -422 -212 -410
rect -246 -444 -212 -422
rect -246 -490 -212 -482
rect -246 -516 -212 -490
rect 212 428 246 454
rect 212 420 246 428
rect 212 360 246 382
rect 212 348 246 360
rect 212 292 246 310
rect 212 276 246 292
rect 212 224 246 238
rect 212 204 246 224
rect 212 156 246 166
rect 212 132 246 156
rect 212 88 246 94
rect 212 60 246 88
rect 212 20 246 22
rect 212 -12 246 20
rect 212 -82 246 -50
rect 212 -84 246 -82
rect 212 -150 246 -122
rect 212 -156 246 -150
rect 212 -218 246 -194
rect 212 -228 246 -218
rect 212 -286 246 -266
rect 212 -300 246 -286
rect 212 -354 246 -338
rect 212 -372 246 -354
rect 212 -422 246 -410
rect 212 -444 246 -422
rect 212 -490 246 -482
rect 212 -516 246 -490
<< metal1 >>
rect -196 541 196 547
rect -196 507 -161 541
rect -127 507 -89 541
rect -55 507 -17 541
rect 17 507 55 541
rect 89 507 127 541
rect 161 507 196 541
rect -196 501 196 507
rect -252 454 -206 469
rect -252 420 -246 454
rect -212 420 -206 454
rect -252 382 -206 420
rect -252 348 -246 382
rect -212 348 -206 382
rect -252 310 -206 348
rect -252 276 -246 310
rect -212 276 -206 310
rect -252 238 -206 276
rect -252 204 -246 238
rect -212 204 -206 238
rect -252 166 -206 204
rect -252 132 -246 166
rect -212 132 -206 166
rect -252 94 -206 132
rect -252 60 -246 94
rect -212 60 -206 94
rect -252 22 -206 60
rect -252 -12 -246 22
rect -212 -12 -206 22
rect -252 -50 -206 -12
rect -252 -84 -246 -50
rect -212 -84 -206 -50
rect -252 -122 -206 -84
rect -252 -156 -246 -122
rect -212 -156 -206 -122
rect -252 -194 -206 -156
rect -252 -228 -246 -194
rect -212 -228 -206 -194
rect -252 -266 -206 -228
rect -252 -300 -246 -266
rect -212 -300 -206 -266
rect -252 -338 -206 -300
rect -252 -372 -246 -338
rect -212 -372 -206 -338
rect -252 -410 -206 -372
rect -252 -444 -246 -410
rect -212 -444 -206 -410
rect -252 -482 -206 -444
rect -252 -516 -246 -482
rect -212 -516 -206 -482
rect -252 -531 -206 -516
rect 206 454 252 469
rect 206 420 212 454
rect 246 420 252 454
rect 206 382 252 420
rect 206 348 212 382
rect 246 348 252 382
rect 206 310 252 348
rect 206 276 212 310
rect 246 276 252 310
rect 206 238 252 276
rect 206 204 212 238
rect 246 204 252 238
rect 206 166 252 204
rect 206 132 212 166
rect 246 132 252 166
rect 206 94 252 132
rect 206 60 212 94
rect 246 60 252 94
rect 206 22 252 60
rect 206 -12 212 22
rect 246 -12 252 22
rect 206 -50 252 -12
rect 206 -84 212 -50
rect 246 -84 252 -50
rect 206 -122 252 -84
rect 206 -156 212 -122
rect 246 -156 252 -122
rect 206 -194 252 -156
rect 206 -228 212 -194
rect 246 -228 252 -194
rect 206 -266 252 -228
rect 206 -300 212 -266
rect 246 -300 252 -266
rect 206 -338 252 -300
rect 206 -372 212 -338
rect 246 -372 252 -338
rect 206 -410 252 -372
rect 206 -444 212 -410
rect 246 -444 252 -410
rect 206 -482 252 -444
rect 206 -516 212 -482
rect 246 -516 252 -482
rect 206 -531 252 -516
<< properties >>
string FIXED_BBOX -343 -626 343 626
<< end >>
