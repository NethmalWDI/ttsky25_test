magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -1094 -198 1094 164
<< pmoslvt >>
rect -1000 -136 1000 64
<< pdiff >>
rect -1058 15 -1000 64
rect -1058 -19 -1046 15
rect -1012 -19 -1000 15
rect -1058 -53 -1000 -19
rect -1058 -87 -1046 -53
rect -1012 -87 -1000 -53
rect -1058 -136 -1000 -87
rect 1000 15 1058 64
rect 1000 -19 1012 15
rect 1046 -19 1058 15
rect 1000 -53 1058 -19
rect 1000 -87 1012 -53
rect 1046 -87 1058 -53
rect 1000 -136 1058 -87
<< pdiffc >>
rect -1046 -19 -1012 15
rect -1046 -87 -1012 -53
rect 1012 -19 1046 15
rect 1012 -87 1046 -53
<< poly >>
rect -705 145 705 161
rect -705 128 -663 145
rect -1000 111 -663 128
rect -629 111 -595 145
rect -561 111 -527 145
rect -493 111 -459 145
rect -425 111 -391 145
rect -357 111 -323 145
rect -289 111 -255 145
rect -221 111 -187 145
rect -153 111 -119 145
rect -85 111 -51 145
rect -17 111 17 145
rect 51 111 85 145
rect 119 111 153 145
rect 187 111 221 145
rect 255 111 289 145
rect 323 111 357 145
rect 391 111 425 145
rect 459 111 493 145
rect 527 111 561 145
rect 595 111 629 145
rect 663 128 705 145
rect 663 111 1000 128
rect -1000 64 1000 111
rect -1000 -162 1000 -136
<< polycont >>
rect -663 111 -629 145
rect -595 111 -561 145
rect -527 111 -493 145
rect -459 111 -425 145
rect -391 111 -357 145
rect -323 111 -289 145
rect -255 111 -221 145
rect -187 111 -153 145
rect -119 111 -85 145
rect -51 111 -17 145
rect 17 111 51 145
rect 85 111 119 145
rect 153 111 187 145
rect 221 111 255 145
rect 289 111 323 145
rect 357 111 391 145
rect 425 111 459 145
rect 493 111 527 145
rect 561 111 595 145
rect 629 111 663 145
<< locali >>
rect -705 111 -665 145
rect -629 111 -595 145
rect -559 111 -527 145
rect -487 111 -459 145
rect -415 111 -391 145
rect -343 111 -323 145
rect -271 111 -255 145
rect -199 111 -187 145
rect -127 111 -119 145
rect -55 111 -51 145
rect 51 111 55 145
rect 119 111 127 145
rect 187 111 199 145
rect 255 111 271 145
rect 323 111 343 145
rect 391 111 415 145
rect 459 111 487 145
rect 527 111 559 145
rect 595 111 629 145
rect 665 111 705 145
rect -1046 17 -1012 42
rect -1046 -53 -1012 -19
rect -1046 -114 -1012 -89
rect 1012 17 1046 42
rect 1012 -53 1046 -19
rect 1012 -114 1046 -89
<< viali >>
rect -665 111 -663 145
rect -663 111 -631 145
rect -593 111 -561 145
rect -561 111 -559 145
rect -521 111 -493 145
rect -493 111 -487 145
rect -449 111 -425 145
rect -425 111 -415 145
rect -377 111 -357 145
rect -357 111 -343 145
rect -305 111 -289 145
rect -289 111 -271 145
rect -233 111 -221 145
rect -221 111 -199 145
rect -161 111 -153 145
rect -153 111 -127 145
rect -89 111 -85 145
rect -85 111 -55 145
rect -17 111 17 145
rect 55 111 85 145
rect 85 111 89 145
rect 127 111 153 145
rect 153 111 161 145
rect 199 111 221 145
rect 221 111 233 145
rect 271 111 289 145
rect 289 111 305 145
rect 343 111 357 145
rect 357 111 377 145
rect 415 111 425 145
rect 425 111 449 145
rect 487 111 493 145
rect 493 111 521 145
rect 559 111 561 145
rect 561 111 593 145
rect 631 111 663 145
rect 663 111 665 145
rect -1046 15 -1012 17
rect -1046 -17 -1012 15
rect -1046 -87 -1012 -55
rect -1046 -89 -1012 -87
rect 1012 15 1046 17
rect 1012 -17 1046 15
rect 1012 -87 1046 -55
rect 1012 -89 1046 -87
<< metal1 >>
rect -701 145 701 151
rect -701 111 -665 145
rect -631 111 -593 145
rect -559 111 -521 145
rect -487 111 -449 145
rect -415 111 -377 145
rect -343 111 -305 145
rect -271 111 -233 145
rect -199 111 -161 145
rect -127 111 -89 145
rect -55 111 -17 145
rect 17 111 55 145
rect 89 111 127 145
rect 161 111 199 145
rect 233 111 271 145
rect 305 111 343 145
rect 377 111 415 145
rect 449 111 487 145
rect 521 111 559 145
rect 593 111 631 145
rect 665 111 701 145
rect -701 105 701 111
rect -1052 17 -1006 38
rect -1052 -17 -1046 17
rect -1012 -17 -1006 17
rect -1052 -55 -1006 -17
rect -1052 -89 -1046 -55
rect -1012 -89 -1006 -55
rect -1052 -110 -1006 -89
rect 1006 17 1052 38
rect 1006 -17 1012 17
rect 1046 -17 1052 17
rect 1006 -55 1052 -17
rect 1006 -89 1012 -55
rect 1046 -89 1052 -55
rect 1006 -110 1052 -89
<< end >>
