magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -396 -384 396 384
<< pmoslvt >>
rect -200 -236 200 164
<< pdiff >>
rect -258 151 -200 164
rect -258 117 -246 151
rect -212 117 -200 151
rect -258 83 -200 117
rect -258 49 -246 83
rect -212 49 -200 83
rect -258 15 -200 49
rect -258 -19 -246 15
rect -212 -19 -200 15
rect -258 -53 -200 -19
rect -258 -87 -246 -53
rect -212 -87 -200 -53
rect -258 -121 -200 -87
rect -258 -155 -246 -121
rect -212 -155 -200 -121
rect -258 -189 -200 -155
rect -258 -223 -246 -189
rect -212 -223 -200 -189
rect -258 -236 -200 -223
rect 200 151 258 164
rect 200 117 212 151
rect 246 117 258 151
rect 200 83 258 117
rect 200 49 212 83
rect 246 49 258 83
rect 200 15 258 49
rect 200 -19 212 15
rect 246 -19 258 15
rect 200 -53 258 -19
rect 200 -87 212 -53
rect 246 -87 258 -53
rect 200 -121 258 -87
rect 200 -155 212 -121
rect 246 -155 258 -121
rect 200 -189 258 -155
rect 200 -223 212 -189
rect 246 -223 258 -189
rect 200 -236 258 -223
<< pdiffc >>
rect -246 117 -212 151
rect -246 49 -212 83
rect -246 -19 -212 15
rect -246 -87 -212 -53
rect -246 -155 -212 -121
rect -246 -223 -212 -189
rect 212 117 246 151
rect 212 49 246 83
rect 212 -19 246 15
rect 212 -87 246 -53
rect 212 -155 246 -121
rect 212 -223 246 -189
<< nsubdiff >>
rect -360 314 360 348
rect -360 221 -326 314
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect -360 -314 -326 -221
rect 326 -314 360 314
rect -360 -348 360 -314
<< nsubdiffcont >>
rect -360 187 -326 221
rect -360 119 -326 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -360 -153 -326 -119
rect -360 -221 -326 -187
<< poly >>
rect -200 245 200 261
rect -200 211 -153 245
rect -119 211 -85 245
rect -51 211 -17 245
rect 17 211 51 245
rect 85 211 119 245
rect 153 211 200 245
rect -200 164 200 211
rect -200 -262 200 -236
<< polycont >>
rect -153 211 -119 245
rect -85 211 -51 245
rect -17 211 17 245
rect 51 211 85 245
rect 119 211 153 245
<< locali >>
rect -360 314 360 348
rect -360 221 -326 314
rect -200 211 -161 245
rect -119 211 -89 245
rect -51 211 -17 245
rect 17 211 51 245
rect 89 211 119 245
rect 161 211 200 245
rect -360 153 -326 187
rect -360 85 -326 119
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect -360 -187 -326 -153
rect -360 -314 -326 -221
rect -246 151 -212 168
rect -246 83 -212 91
rect -246 15 -212 19
rect -246 -91 -212 -87
rect -246 -163 -212 -155
rect -246 -240 -212 -223
rect 212 151 246 168
rect 212 83 246 91
rect 212 15 246 19
rect 212 -91 246 -87
rect 212 -163 246 -155
rect 212 -240 246 -223
rect 326 -314 360 314
rect -360 -348 360 -314
<< viali >>
rect -161 211 -153 245
rect -153 211 -127 245
rect -89 211 -85 245
rect -85 211 -55 245
rect -17 211 17 245
rect 55 211 85 245
rect 85 211 89 245
rect 127 211 153 245
rect 153 211 161 245
rect -246 117 -212 125
rect -246 91 -212 117
rect -246 49 -212 53
rect -246 19 -212 49
rect -246 -53 -212 -19
rect -246 -121 -212 -91
rect -246 -125 -212 -121
rect -246 -189 -212 -163
rect -246 -197 -212 -189
rect 212 117 246 125
rect 212 91 246 117
rect 212 49 246 53
rect 212 19 246 49
rect 212 -53 246 -19
rect 212 -121 246 -91
rect 212 -125 246 -121
rect 212 -189 246 -163
rect 212 -197 246 -189
<< metal1 >>
rect -196 245 196 251
rect -196 211 -161 245
rect -127 211 -89 245
rect -55 211 -17 245
rect 17 211 55 245
rect 89 211 127 245
rect 161 211 196 245
rect -196 205 196 211
rect -252 125 -206 164
rect -252 91 -246 125
rect -212 91 -206 125
rect -252 53 -206 91
rect -252 19 -246 53
rect -212 19 -206 53
rect -252 -19 -206 19
rect -252 -53 -246 -19
rect -212 -53 -206 -19
rect -252 -91 -206 -53
rect -252 -125 -246 -91
rect -212 -125 -206 -91
rect -252 -163 -206 -125
rect -252 -197 -246 -163
rect -212 -197 -206 -163
rect -252 -236 -206 -197
rect 206 125 252 164
rect 206 91 212 125
rect 246 91 252 125
rect 206 53 252 91
rect 206 19 212 53
rect 246 19 252 53
rect 206 -19 252 19
rect 206 -53 212 -19
rect 246 -53 252 -19
rect 206 -91 252 -53
rect 206 -125 212 -91
rect 246 -125 252 -91
rect 206 -163 252 -125
rect 206 -197 212 -163
rect 246 -197 252 -163
rect 206 -236 252 -197
<< properties >>
string FIXED_BBOX -343 -331 343 331
<< end >>
