magic
tech sky130A
magscale 1 2
timestamp 1757164387
<< metal2 >>
rect 27170 45058 27270 45080
rect 27170 45002 27192 45058
rect 27248 45002 27270 45058
rect 27170 44980 27270 45002
rect 27720 45058 27820 45080
rect 27720 45002 27742 45058
rect 27798 45002 27820 45058
rect 27720 44980 27820 45002
rect 27210 44830 27270 44980
rect 27760 44930 27820 44980
rect 27760 44903 29810 44930
rect 27760 44870 29712 44903
rect 29670 44847 29712 44870
rect 29768 44847 29810 44903
rect 29670 44830 29810 44847
rect 27210 44780 29610 44830
rect 29470 44753 29610 44780
rect 29470 44697 29512 44753
rect 29568 44697 29610 44753
rect 29470 44680 29610 44697
<< via2 >>
rect 27192 45002 27248 45058
rect 27742 45002 27798 45058
rect 29712 44847 29768 44903
rect 29512 44697 29568 44753
<< metal3 >>
rect 27170 45062 27270 45080
rect 27170 44998 27188 45062
rect 27252 44998 27270 45062
rect 27170 44980 27270 44998
rect 27720 45062 27820 45080
rect 27720 44998 27738 45062
rect 27802 44998 27820 45062
rect 27720 44980 27820 44998
rect 29670 44907 29810 44930
rect 29670 44903 29713 44907
rect 29670 44847 29712 44903
rect 29670 44843 29713 44847
rect 29777 44843 29810 44907
rect 29670 44830 29810 44843
rect 29470 44757 29610 44770
rect 29470 44693 29508 44757
rect 29572 44693 29610 44757
rect 29470 44680 29610 44693
rect 200 13572 4770 13620
rect 200 13508 253 13572
rect 317 13508 433 13572
rect 497 13508 4770 13572
rect 200 13432 4770 13508
rect 200 13368 253 13432
rect 317 13368 433 13432
rect 497 13368 4770 13432
rect 200 13320 4770 13368
rect 27980 7930 28300 8010
rect 27980 7892 29610 7930
rect 27980 7828 29508 7892
rect 29572 7828 29610 7892
rect 27980 7790 29610 7828
rect 27980 7710 28300 7790
rect 27970 7472 29810 7510
rect 27970 7408 29708 7472
rect 29772 7408 29810 7472
rect 27970 7370 29810 7408
rect 27970 7210 28280 7370
rect 200 3157 3940 3190
rect 200 3093 243 3157
rect 307 3093 373 3157
rect 437 3093 503 3157
rect 567 3142 3940 3157
rect 567 3093 3678 3142
rect 200 3078 3678 3093
rect 3742 3078 3828 3142
rect 3892 3078 3940 3142
rect 200 3002 3940 3078
rect 200 2997 3678 3002
rect 200 2933 243 2997
rect 307 2933 373 2997
rect 437 2933 503 2997
rect 567 2938 3678 2997
rect 3742 2938 3828 3002
rect 3892 2938 3940 3002
rect 567 2933 3940 2938
rect 200 2890 3940 2933
rect 800 2637 28830 2680
rect 800 2573 833 2637
rect 897 2573 963 2637
rect 1027 2573 1093 2637
rect 1157 2602 28830 2637
rect 1157 2573 28558 2602
rect 800 2538 28558 2573
rect 28622 2538 28708 2602
rect 28772 2538 28830 2602
rect 800 2477 28830 2538
rect 800 2413 833 2477
rect 897 2413 963 2477
rect 1027 2413 1093 2477
rect 1157 2472 28830 2477
rect 1157 2413 28558 2472
rect 800 2408 28558 2413
rect 28622 2408 28708 2472
rect 28772 2408 28830 2472
rect 800 2370 28830 2408
<< via3 >>
rect 27188 45058 27252 45062
rect 27188 45002 27192 45058
rect 27192 45002 27248 45058
rect 27248 45002 27252 45058
rect 27188 44998 27252 45002
rect 27738 45058 27802 45062
rect 27738 45002 27742 45058
rect 27742 45002 27798 45058
rect 27798 45002 27802 45058
rect 27738 44998 27802 45002
rect 29713 44903 29777 44907
rect 29713 44847 29768 44903
rect 29768 44847 29777 44903
rect 29713 44843 29777 44847
rect 29508 44753 29572 44757
rect 29508 44697 29512 44753
rect 29512 44697 29568 44753
rect 29568 44697 29572 44753
rect 29508 44693 29572 44697
rect 253 13508 317 13572
rect 433 13508 497 13572
rect 253 13368 317 13432
rect 433 13368 497 13432
rect 29508 7828 29572 7892
rect 29708 7408 29772 7472
rect 243 3093 307 3157
rect 373 3093 437 3157
rect 503 3093 567 3157
rect 3678 3078 3742 3142
rect 3828 3078 3892 3142
rect 243 2933 307 2997
rect 373 2933 437 2997
rect 503 2933 567 2997
rect 3678 2938 3742 3002
rect 3828 2938 3892 3002
rect 833 2573 897 2637
rect 963 2573 1027 2637
rect 1093 2573 1157 2637
rect 28558 2538 28622 2602
rect 28708 2538 28772 2602
rect 833 2413 897 2477
rect 963 2413 1027 2477
rect 1093 2413 1157 2477
rect 28558 2408 28622 2472
rect 28708 2408 28772 2472
<< metal4 >>
rect 6134 44810 6194 45152
rect 6686 44810 6746 45152
rect 7238 44810 7298 45152
rect 7790 44810 7850 45152
rect 8342 44810 8402 45152
rect 8894 44810 8954 45152
rect 9446 44810 9506 45152
rect 9998 44810 10058 45152
rect 10550 44810 10610 45152
rect 11102 44810 11162 45152
rect 11654 44810 11714 45152
rect 12206 44810 12266 45152
rect 12758 44810 12818 45152
rect 13310 44810 13370 45152
rect 13862 44810 13922 45152
rect 14414 45040 14474 45152
rect 14966 45040 15026 45152
rect 15518 45040 15578 45152
rect 16070 45040 16130 45152
rect 16622 45040 16682 45152
rect 17174 45040 17234 45152
rect 17726 45040 17786 45152
rect 18278 45040 18338 45152
rect 18830 45040 18890 45152
rect 19382 45040 19442 45152
rect 19934 45040 19994 45152
rect 20486 45040 20546 45152
rect 21038 45040 21098 45152
rect 21590 45040 21650 45152
rect 22142 45040 22202 45152
rect 22694 45040 22754 45152
rect 23246 45040 23306 45152
rect 23798 45040 23858 45152
rect 24350 45040 24410 45152
rect 24902 45040 24962 45152
rect 25454 45040 25514 45152
rect 26006 45040 26066 45152
rect 26558 45040 26618 45152
rect 14176 44980 26618 45040
rect 14176 44810 14236 44980
rect 14414 44952 14474 44980
rect 14966 44952 15026 44980
rect 15518 44952 15578 44980
rect 16070 44952 16130 44980
rect 16622 44952 16682 44980
rect 17174 44952 17234 44980
rect 17726 44952 17786 44980
rect 18278 44952 18338 44980
rect 18830 44952 18890 44980
rect 19382 44952 19442 44980
rect 19934 44952 19994 44980
rect 20486 44952 20546 44980
rect 21038 44952 21098 44980
rect 21590 44952 21650 44980
rect 22142 44952 22202 44980
rect 22694 44952 22754 44980
rect 23246 44952 23306 44980
rect 23798 44952 23858 44980
rect 24350 44952 24410 44980
rect 24902 44952 24962 44980
rect 25454 44952 25514 44980
rect 26006 44952 26066 44980
rect 800 44510 14236 44810
rect 26558 44770 26618 44980
rect 27110 45080 27170 45152
rect 27662 45080 27722 45152
rect 27110 45062 27270 45080
rect 27110 44998 27188 45062
rect 27252 44998 27270 45062
rect 27110 44980 27270 44998
rect 27662 45062 27820 45080
rect 27662 44998 27738 45062
rect 27802 44998 27820 45062
rect 27662 44980 27820 44998
rect 28214 45060 28274 45152
rect 28766 45060 28826 45152
rect 29318 45060 29378 45152
rect 28214 45000 29378 45060
rect 27110 44920 27170 44980
rect 27662 44930 27722 44980
rect 28214 44770 28274 45000
rect 28766 44952 28826 45000
rect 29318 44952 29378 45000
rect 29670 44907 29810 44930
rect 29670 44843 29713 44907
rect 29777 44843 29810 44907
rect 26558 44710 28274 44770
rect 29470 44757 29610 44780
rect 200 13572 600 44152
rect 200 13508 253 13572
rect 317 13508 433 13572
rect 497 13508 600 13572
rect 200 13432 600 13508
rect 200 13368 253 13432
rect 317 13368 433 13432
rect 497 13368 600 13432
rect 200 3157 600 13368
rect 200 3093 243 3157
rect 307 3093 373 3157
rect 437 3093 503 3157
rect 567 3093 600 3157
rect 200 2997 600 3093
rect 200 2933 243 2997
rect 307 2933 373 2997
rect 437 2933 503 2997
rect 567 2933 600 2997
rect 200 1000 600 2933
rect 800 2637 1200 44510
rect 800 2573 833 2637
rect 897 2573 963 2637
rect 1027 2573 1093 2637
rect 1157 2573 1200 2637
rect 800 2477 1200 2573
rect 800 2413 833 2477
rect 897 2413 963 2477
rect 1027 2413 1093 2477
rect 1157 2413 1200 2477
rect 800 1000 1200 2413
rect 2650 44150 13386 44450
rect 2650 1401 2950 44150
rect 3050 43770 13006 44070
rect 3050 1977 3350 43770
rect 13936 37550 14236 44510
rect 29470 44693 29508 44757
rect 29572 44693 29610 44757
rect 13936 36930 14236 37430
rect 15080 36470 15210 36570
rect 29470 7892 29610 44693
rect 29470 7828 29508 7892
rect 29572 7828 29610 7892
rect 29470 7790 29610 7828
rect 29670 7472 29810 44843
rect 29670 7408 29708 7472
rect 29772 7408 29810 7472
rect 29670 7370 29810 7408
rect 3660 3142 3760 3160
rect 3660 3078 3678 3142
rect 3742 3078 3760 3142
rect 3660 3060 3760 3078
rect 3810 3142 3910 3160
rect 3810 3078 3828 3142
rect 3892 3078 3910 3142
rect 3810 3060 3910 3078
rect 3660 3002 3760 3020
rect 3660 2938 3678 3002
rect 3742 2938 3760 3002
rect 3660 2920 3760 2938
rect 3810 3002 3910 3020
rect 3810 2938 3828 3002
rect 3892 2938 3910 3002
rect 3810 2920 3910 2938
rect 3050 1677 15084 1977
rect 2650 1101 11220 1401
rect 11040 200 11220 1101
rect 14904 200 15084 1677
rect 17676 1134 17976 3310
rect 18976 1654 19276 3507
rect 19516 2179 19816 3336
rect 28526 2602 28826 3099
rect 28526 2538 28558 2602
rect 28622 2538 28708 2602
rect 28772 2538 28826 2602
rect 28526 2472 28826 2538
rect 28526 2408 28558 2472
rect 28622 2408 28708 2472
rect 28772 2408 28826 2472
rect 28526 2372 28826 2408
rect 19516 1878 26678 2179
rect 18976 1354 22812 1654
rect 17676 834 18950 1134
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11040 0 11222 200
rect 14904 1 15086 200
rect 14906 0 15086 1
rect 18770 0 18950 834
rect 22632 200 22812 1354
rect 22632 0 22814 200
rect 26498 0 26678 1878
rect 29056 1070 29356 3060
rect 29056 770 30542 1070
rect 30362 0 30542 770
use op_amp_lvs_final  op_amp_lvs_final_0 /foss/designs
timestamp 1585778769
transform 0 -1 29156 1 0 2890
box -130 -200 41812 25723
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 600 90 0 0 clk
port 4 nsew
flabel metal4 s 28796 45052 28796 45052 0 FreeSans 600 90 0 0 clk
flabel metal4 s 28796 45052 28796 45052 0 FreeSans 600 90 0 0 clk
flabel metal4 s 28796 45052 28796 45052 0 FreeSans 600 90 0 0 clk
flabel metal4 s 28796 45052 28796 45052 0 FreeSans 600 90 0 0 clk
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 600 90 0 0 ena
port 5 nsew
flabel metal4 s 29348 45052 29348 45052 0 FreeSans 600 90 0 0 ena
flabel metal4 s 29348 45052 29348 45052 0 FreeSans 600 90 0 0 ena
flabel metal4 s 29348 45052 29348 45052 0 FreeSans 600 90 0 0 ena
flabel metal4 s 29348 45052 29348 45052 0 FreeSans 600 90 0 0 ena
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 600 90 0 0 rst_n
port 1 nsew
flabel metal4 s 28244 45052 28244 45052 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 28244 45052 28244 45052 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 28244 45052 28244 45052 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 28244 45052 28244 45052 0 FreeSans 600 90 0 0 rst_n
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 600 90 0 0 ui_in[0]
port 6 nsew
flabel metal4 s 27692 45052 27692 45052 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 27692 45052 27692 45052 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 27692 45052 27692 45052 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 27692 45052 27692 45052 0 FreeSans 600 90 0 0 ui_in[0]
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 600 90 0 0 ui_in[1]
port 7 nsew
flabel metal4 s 27140 45052 27140 45052 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 27140 45052 27140 45052 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 27140 45052 27140 45052 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 27140 45052 27140 45052 0 FreeSans 600 90 0 0 ui_in[1]
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 600 90 0 0 ui_in[2]
port 8 nsew
flabel metal4 s 26588 45052 26588 45052 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 26588 45052 26588 45052 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 26588 45052 26588 45052 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 26588 45052 26588 45052 0 FreeSans 600 90 0 0 ui_in[2]
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 600 90 0 0 ui_in[3]
port 9 nsew
flabel metal4 s 26036 45052 26036 45052 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 26036 45052 26036 45052 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 26036 45052 26036 45052 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 26036 45052 26036 45052 0 FreeSans 600 90 0 0 ui_in[3]
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 600 90 0 0 ui_in[4]
port 10 nsew
flabel metal4 s 25484 45052 25484 45052 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 25484 45052 25484 45052 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 25484 45052 25484 45052 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 25484 45052 25484 45052 0 FreeSans 600 90 0 0 ui_in[4]
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 600 90 0 0 ui_in[5]
port 11 nsew
flabel metal4 s 24932 45052 24932 45052 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 24932 45052 24932 45052 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 24932 45052 24932 45052 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 24932 45052 24932 45052 0 FreeSans 600 90 0 0 ui_in[5]
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 600 90 0 0 ui_in[6]
port 12 nsew
flabel metal4 s 24380 45052 24380 45052 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 24380 45052 24380 45052 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 24380 45052 24380 45052 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 24380 45052 24380 45052 0 FreeSans 600 90 0 0 ui_in[6]
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 600 90 0 0 ui_in[7]
port 13 nsew
flabel metal4 s 23828 45052 23828 45052 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 23828 45052 23828 45052 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 23828 45052 23828 45052 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 23828 45052 23828 45052 0 FreeSans 600 90 0 0 ui_in[7]
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 600 90 0 0 uio_in[0]
port 14 nsew
flabel metal4 s 23276 45052 23276 45052 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 23276 45052 23276 45052 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 23276 45052 23276 45052 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 23276 45052 23276 45052 0 FreeSans 600 90 0 0 uio_in[0]
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 600 90 0 0 uio_in[1]
port 15 nsew
flabel metal4 s 22724 45052 22724 45052 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22724 45052 22724 45052 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22724 45052 22724 45052 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22724 45052 22724 45052 0 FreeSans 600 90 0 0 uio_in[1]
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 600 90 0 0 uio_in[2]
port 16 nsew
flabel metal4 s 22172 45052 22172 45052 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 22172 45052 22172 45052 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 22172 45052 22172 45052 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 22172 45052 22172 45052 0 FreeSans 600 90 0 0 uio_in[2]
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 600 90 0 0 uio_in[3]
port 17 nsew
flabel metal4 s 21620 45052 21620 45052 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 21620 45052 21620 45052 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 21620 45052 21620 45052 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 21620 45052 21620 45052 0 FreeSans 600 90 0 0 uio_in[3]
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 600 90 0 0 uio_in[4]
port 18 nsew
flabel metal4 s 21068 45052 21068 45052 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 21068 45052 21068 45052 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 21068 45052 21068 45052 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 21068 45052 21068 45052 0 FreeSans 600 90 0 0 uio_in[4]
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 600 90 0 0 uio_in[5]
port 19 nsew
flabel metal4 s 20516 45052 20516 45052 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 20516 45052 20516 45052 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 20516 45052 20516 45052 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 20516 45052 20516 45052 0 FreeSans 600 90 0 0 uio_in[5]
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 600 90 0 0 uio_in[6]
port 20 nsew
flabel metal4 s 19964 45052 19964 45052 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 19964 45052 19964 45052 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 19964 45052 19964 45052 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 19964 45052 19964 45052 0 FreeSans 600 90 0 0 uio_in[6]
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 600 90 0 0 uio_in[7]
port 21 nsew
flabel metal4 s 19412 45052 19412 45052 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 19412 45052 19412 45052 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 19412 45052 19412 45052 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 19412 45052 19412 45052 0 FreeSans 600 90 0 0 uio_in[7]
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 600 90 0 0 uo_out[0]
port 22 nsew
flabel metal4 s 18860 45052 18860 45052 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 18860 45052 18860 45052 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 18860 45052 18860 45052 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 18860 45052 18860 45052 0 FreeSans 600 90 0 0 uo_out[0]
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 600 90 0 0 uo_out[1]
port 23 nsew
flabel metal4 s 18308 45052 18308 45052 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 18308 45052 18308 45052 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 18308 45052 18308 45052 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 18308 45052 18308 45052 0 FreeSans 600 90 0 0 uo_out[1]
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 600 90 0 0 uo_out[2]
port 24 nsew
flabel metal4 s 17756 45052 17756 45052 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 17756 45052 17756 45052 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 17756 45052 17756 45052 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 17756 45052 17756 45052 0 FreeSans 600 90 0 0 uo_out[2]
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 600 90 0 0 uo_out[3]
port 25 nsew
flabel metal4 s 17204 45052 17204 45052 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 17204 45052 17204 45052 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 17204 45052 17204 45052 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 17204 45052 17204 45052 0 FreeSans 600 90 0 0 uo_out[3]
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 600 90 0 0 uo_out[4]
port 26 nsew
flabel metal4 s 16652 45052 16652 45052 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 16652 45052 16652 45052 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 16652 45052 16652 45052 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 16652 45052 16652 45052 0 FreeSans 600 90 0 0 uo_out[4]
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 600 90 0 0 uo_out[5]
port 27 nsew
flabel metal4 s 16100 45052 16100 45052 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 16100 45052 16100 45052 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 16100 45052 16100 45052 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 16100 45052 16100 45052 0 FreeSans 600 90 0 0 uo_out[5]
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 600 90 0 0 uo_out[6]
port 28 nsew
flabel metal4 s 15548 45052 15548 45052 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 15548 45052 15548 45052 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 15548 45052 15548 45052 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 15548 45052 15548 45052 0 FreeSans 600 90 0 0 uo_out[6]
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 600 90 0 0 uio_oe[7]
port 29 nsew
flabel metal4 s 6164 45052 6164 45052 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 6164 45052 6164 45052 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 6164 45052 6164 45052 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 6164 45052 6164 45052 0 FreeSans 600 90 0 0 uio_oe[7]
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 600 90 0 0 uio_out[0]
port 30 nsew
flabel metal4 s 14444 45052 14444 45052 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 14444 45052 14444 45052 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 14444 45052 14444 45052 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 14444 45052 14444 45052 0 FreeSans 600 90 0 0 uio_out[0]
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 600 90 0 0 uio_out[1]
port 31 nsew
flabel metal4 s 13892 45052 13892 45052 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 13892 45052 13892 45052 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 13892 45052 13892 45052 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 13892 45052 13892 45052 0 FreeSans 600 90 0 0 uio_out[1]
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 600 90 0 0 uio_out[2]
port 32 nsew
flabel metal4 s 13340 45052 13340 45052 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 13340 45052 13340 45052 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 13340 45052 13340 45052 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 13340 45052 13340 45052 0 FreeSans 600 90 0 0 uio_out[2]
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 600 90 0 0 uio_out[3]
port 33 nsew
flabel metal4 s 12788 45052 12788 45052 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 12788 45052 12788 45052 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 12788 45052 12788 45052 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 12788 45052 12788 45052 0 FreeSans 600 90 0 0 uio_out[3]
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 600 90 0 0 uio_out[4]
port 34 nsew
flabel metal4 s 12236 45052 12236 45052 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 12236 45052 12236 45052 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 12236 45052 12236 45052 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 12236 45052 12236 45052 0 FreeSans 600 90 0 0 uio_out[4]
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 600 90 0 0 uio_out[5]
port 35 nsew
flabel metal4 s 11684 45052 11684 45052 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 11684 45052 11684 45052 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 11684 45052 11684 45052 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 11684 45052 11684 45052 0 FreeSans 600 90 0 0 uio_out[5]
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 600 90 0 0 uio_out[6]
port 36 nsew
flabel metal4 s 11132 45052 11132 45052 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 11132 45052 11132 45052 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 11132 45052 11132 45052 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 11132 45052 11132 45052 0 FreeSans 600 90 0 0 uio_out[6]
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 600 90 0 0 uio_out[7]
port 37 nsew
flabel metal4 s 10580 45052 10580 45052 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 10580 45052 10580 45052 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 10580 45052 10580 45052 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 10580 45052 10580 45052 0 FreeSans 600 90 0 0 uio_out[7]
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 600 90 0 0 uio_oe[0]
port 38 nsew
flabel metal4 s 10028 45052 10028 45052 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 10028 45052 10028 45052 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 10028 45052 10028 45052 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 10028 45052 10028 45052 0 FreeSans 600 90 0 0 uio_oe[0]
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 600 90 0 0 uio_oe[1]
port 39 nsew
flabel metal4 s 9476 45052 9476 45052 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 9476 45052 9476 45052 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 9476 45052 9476 45052 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 9476 45052 9476 45052 0 FreeSans 600 90 0 0 uio_oe[1]
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 600 90 0 0 uio_oe[2]
port 40 nsew
flabel metal4 s 8924 45052 8924 45052 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 8924 45052 8924 45052 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 8924 45052 8924 45052 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 8924 45052 8924 45052 0 FreeSans 600 90 0 0 uio_oe[2]
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 600 90 0 0 uio_oe[3]
port 41 nsew
flabel metal4 s 8372 45052 8372 45052 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 8372 45052 8372 45052 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 8372 45052 8372 45052 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 8372 45052 8372 45052 0 FreeSans 600 90 0 0 uio_oe[3]
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 600 90 0 0 uio_oe[4]
port 42 nsew
flabel metal4 s 7820 45052 7820 45052 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 7820 45052 7820 45052 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 7820 45052 7820 45052 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 7820 45052 7820 45052 0 FreeSans 600 90 0 0 uio_oe[4]
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 600 90 0 0 uio_oe[5]
port 43 nsew
flabel metal4 s 7268 45052 7268 45052 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 7268 45052 7268 45052 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 7268 45052 7268 45052 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 7268 45052 7268 45052 0 FreeSans 600 90 0 0 uio_oe[5]
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 600 90 0 0 uio_oe[6]
port 44 nsew
flabel metal4 s 6716 45052 6716 45052 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 6716 45052 6716 45052 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 6716 45052 6716 45052 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 6716 45052 6716 45052 0 FreeSans 600 90 0 0 uio_oe[6]
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 600 90 0 0 uo_out[7]
port 45 nsew
flabel metal4 s 14996 45052 14996 45052 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 14996 45052 14996 45052 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 14996 45052 14996 45052 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 14996 45052 14996 45052 0 FreeSans 600 90 0 0 uo_out[7]
flabel metal4 s 14906 0 15086 200 0 FreeSans 1200 0 0 0 ua[4]
port 46 nsew
flabel metal4 s 14996 100 14996 100 0 FreeSans 1200 0 0 0 ua[4]
flabel metal4 s 14996 100 14996 100 0 FreeSans 1200 0 0 0 ua[4]
flabel metal4 s 14996 100 14996 100 0 FreeSans 1200 0 0 0 ua[4]
flabel metal4 s 14996 100 14996 100 0 FreeSans 1200 0 0 0 ua[4]
flabel metal4 s 11042 0 11222 200 0 FreeSans 1200 0 0 0 ua[5]
port 47 nsew
flabel metal4 s 11132 100 11132 100 0 FreeSans 1200 0 0 0 ua[5]
flabel metal4 s 11132 100 11132 100 0 FreeSans 1200 0 0 0 ua[5]
flabel metal4 s 11132 100 11132 100 0 FreeSans 1200 0 0 0 ua[5]
flabel metal4 s 11132 100 11132 100 0 FreeSans 1200 0 0 0 ua[5]
flabel metal4 s 7178 0 7358 200 0 FreeSans 1200 0 0 0 ua[6]
port 48 nsew
flabel metal4 s 7268 100 7268 100 0 FreeSans 1200 0 0 0 ua[6]
flabel metal4 s 7268 100 7268 100 0 FreeSans 1200 0 0 0 ua[6]
flabel metal4 s 7268 100 7268 100 0 FreeSans 1200 0 0 0 ua[6]
flabel metal4 s 7268 100 7268 100 0 FreeSans 1200 0 0 0 ua[6]
flabel metal4 s 3314 0 3494 200 0 FreeSans 1200 0 0 0 ua[7]
port 49 nsew
flabel metal4 s 3404 100 3404 100 0 FreeSans 1200 0 0 0 ua[7]
flabel metal4 s 3404 100 3404 100 0 FreeSans 1200 0 0 0 ua[7]
flabel metal4 s 3404 100 3404 100 0 FreeSans 1200 0 0 0 ua[7]
flabel metal4 s 3404 100 3404 100 0 FreeSans 1200 0 0 0 ua[7]
flabel metal4 s 200 1000 600 44152 1 FreeSans 500 0 0 0 VDPWR
port 2 nsew
flabel metal4 s 800 1000 1200 44152 1 FreeSans 500 0 0 0 VGND
port 3 nsew
flabel metal4 s 800 1000 1200 1280 0 FreeSans 600 0 0 0 VGND
port 3 nsew
flabel metal4 s 200 1000 600 1220 0 FreeSans 600 0 0 0 VDPWR
port 2 nsew
flabel metal4 s 30362 0 30542 200 0 FreeSans 1200 0 0 0 ua[0]
port 50 nsew
flabel metal4 s 26498 0 26678 200 0 FreeSans 1200 0 0 0 ua[1]
port 51 nsew
flabel metal4 s 26588 100 26588 100 0 FreeSans 1200 0 0 0 ua[1]
flabel metal4 s 26588 100 26588 100 0 FreeSans 1200 0 0 0 ua[1]
flabel metal4 s 26588 100 26588 100 0 FreeSans 1200 0 0 0 ua[1]
flabel metal4 s 26588 100 26588 100 0 FreeSans 1200 0 0 0 ua[1]
flabel metal4 s 22634 0 22814 200 0 FreeSans 1200 0 0 0 ua[2]
port 52 nsew
flabel metal4 s 22724 100 22724 100 0 FreeSans 1200 0 0 0 ua[2]
flabel metal4 s 22724 100 22724 100 0 FreeSans 1200 0 0 0 ua[2]
flabel metal4 s 22724 100 22724 100 0 FreeSans 1200 0 0 0 ua[2]
flabel metal4 s 22724 100 22724 100 0 FreeSans 1200 0 0 0 ua[2]
flabel metal4 s 18770 0 18950 200 0 FreeSans 1200 0 0 0 ua[3]
port 53 nsew
flabel metal4 s 18860 100 18860 100 0 FreeSans 1200 0 0 0 ua[3]
flabel metal4 s 18860 100 18860 100 0 FreeSans 1200 0 0 0 ua[3]
flabel metal4 s 18860 100 18860 100 0 FreeSans 1200 0 0 0 ua[3]
flabel metal4 s 18860 100 18860 100 0 FreeSans 1200 0 0 0 ua[3]
flabel metal4 s 30452 100 30452 100 0 FreeSans 1200 0 0 0 ua[0]
flabel metal4 s 30452 100 30452 100 0 FreeSans 1200 0 0 0 ua[0]
flabel metal4 s 30452 100 30452 100 0 FreeSans 1200 0 0 0 ua[0]
flabel metal4 s 30452 100 30452 100 0 FreeSans 1200 0 0 0 ua[0]
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
