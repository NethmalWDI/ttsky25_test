magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< nwell >>
rect -2196 -284 2196 284
<< pmoslvt >>
rect -2000 -64 2000 136
<< pdiff >>
rect -2058 121 -2000 136
rect -2058 87 -2046 121
rect -2012 87 -2000 121
rect -2058 53 -2000 87
rect -2058 19 -2046 53
rect -2012 19 -2000 53
rect -2058 -15 -2000 19
rect -2058 -49 -2046 -15
rect -2012 -49 -2000 -15
rect -2058 -64 -2000 -49
rect 2000 121 2058 136
rect 2000 87 2012 121
rect 2046 87 2058 121
rect 2000 53 2058 87
rect 2000 19 2012 53
rect 2046 19 2058 53
rect 2000 -15 2058 19
rect 2000 -49 2012 -15
rect 2046 -49 2058 -15
rect 2000 -64 2058 -49
<< pdiffc >>
rect -2046 87 -2012 121
rect -2046 19 -2012 53
rect -2046 -49 -2012 -15
rect 2012 87 2046 121
rect 2012 19 2046 53
rect 2012 -49 2046 -15
<< nsubdiff >>
rect -2160 214 -2057 248
rect -2023 214 -1989 248
rect -1955 214 -1921 248
rect -1887 214 -1853 248
rect -1819 214 -1785 248
rect -1751 214 -1717 248
rect -1683 214 -1649 248
rect -1615 214 -1581 248
rect -1547 214 -1513 248
rect -1479 214 -1445 248
rect -1411 214 -1377 248
rect -1343 214 -1309 248
rect -1275 214 -1241 248
rect -1207 214 -1173 248
rect -1139 214 -1105 248
rect -1071 214 -1037 248
rect -1003 214 -969 248
rect -935 214 -901 248
rect -867 214 -833 248
rect -799 214 -765 248
rect -731 214 -697 248
rect -663 214 -629 248
rect -595 214 -561 248
rect -527 214 -493 248
rect -459 214 -425 248
rect -391 214 -357 248
rect -323 214 -289 248
rect -255 214 -221 248
rect -187 214 -153 248
rect -119 214 -85 248
rect -51 214 -17 248
rect 17 214 51 248
rect 85 214 119 248
rect 153 214 187 248
rect 221 214 255 248
rect 289 214 323 248
rect 357 214 391 248
rect 425 214 459 248
rect 493 214 527 248
rect 561 214 595 248
rect 629 214 663 248
rect 697 214 731 248
rect 765 214 799 248
rect 833 214 867 248
rect 901 214 935 248
rect 969 214 1003 248
rect 1037 214 1071 248
rect 1105 214 1139 248
rect 1173 214 1207 248
rect 1241 214 1275 248
rect 1309 214 1343 248
rect 1377 214 1411 248
rect 1445 214 1479 248
rect 1513 214 1547 248
rect 1581 214 1615 248
rect 1649 214 1683 248
rect 1717 214 1751 248
rect 1785 214 1819 248
rect 1853 214 1887 248
rect 1921 214 1955 248
rect 1989 214 2023 248
rect 2057 214 2160 248
rect -2160 -214 -2126 214
rect 2126 -214 2160 214
rect -2160 -248 2160 -214
<< nsubdiffcont >>
rect -2057 214 -2023 248
rect -1989 214 -1955 248
rect -1921 214 -1887 248
rect -1853 214 -1819 248
rect -1785 214 -1751 248
rect -1717 214 -1683 248
rect -1649 214 -1615 248
rect -1581 214 -1547 248
rect -1513 214 -1479 248
rect -1445 214 -1411 248
rect -1377 214 -1343 248
rect -1309 214 -1275 248
rect -1241 214 -1207 248
rect -1173 214 -1139 248
rect -1105 214 -1071 248
rect -1037 214 -1003 248
rect -969 214 -935 248
rect -901 214 -867 248
rect -833 214 -799 248
rect -765 214 -731 248
rect -697 214 -663 248
rect -629 214 -595 248
rect -561 214 -527 248
rect -493 214 -459 248
rect -425 214 -391 248
rect -357 214 -323 248
rect -289 214 -255 248
rect -221 214 -187 248
rect -153 214 -119 248
rect -85 214 -51 248
rect -17 214 17 248
rect 51 214 85 248
rect 119 214 153 248
rect 187 214 221 248
rect 255 214 289 248
rect 323 214 357 248
rect 391 214 425 248
rect 459 214 493 248
rect 527 214 561 248
rect 595 214 629 248
rect 663 214 697 248
rect 731 214 765 248
rect 799 214 833 248
rect 867 214 901 248
rect 935 214 969 248
rect 1003 214 1037 248
rect 1071 214 1105 248
rect 1139 214 1173 248
rect 1207 214 1241 248
rect 1275 214 1309 248
rect 1343 214 1377 248
rect 1411 214 1445 248
rect 1479 214 1513 248
rect 1547 214 1581 248
rect 1615 214 1649 248
rect 1683 214 1717 248
rect 1751 214 1785 248
rect 1819 214 1853 248
rect 1887 214 1921 248
rect 1955 214 1989 248
rect 2023 214 2057 248
<< poly >>
rect -2000 136 2000 162
rect -2000 -111 2000 -64
rect -2000 -145 -1955 -111
rect -1921 -145 -1887 -111
rect -1853 -145 -1819 -111
rect -1785 -145 -1751 -111
rect -1717 -145 -1683 -111
rect -1649 -145 -1615 -111
rect -1581 -145 -1547 -111
rect -1513 -145 -1479 -111
rect -1445 -145 -1411 -111
rect -1377 -145 -1343 -111
rect -1309 -145 -1275 -111
rect -1241 -145 -1207 -111
rect -1173 -145 -1139 -111
rect -1105 -145 -1071 -111
rect -1037 -145 -1003 -111
rect -969 -145 -935 -111
rect -901 -145 -867 -111
rect -833 -145 -799 -111
rect -765 -145 -731 -111
rect -697 -145 -663 -111
rect -629 -145 -595 -111
rect -561 -145 -527 -111
rect -493 -145 -459 -111
rect -425 -145 -391 -111
rect -357 -145 -323 -111
rect -289 -145 -255 -111
rect -221 -145 -187 -111
rect -153 -145 -119 -111
rect -85 -145 -51 -111
rect -17 -145 17 -111
rect 51 -145 85 -111
rect 119 -145 153 -111
rect 187 -145 221 -111
rect 255 -145 289 -111
rect 323 -145 357 -111
rect 391 -145 425 -111
rect 459 -145 493 -111
rect 527 -145 561 -111
rect 595 -145 629 -111
rect 663 -145 697 -111
rect 731 -145 765 -111
rect 799 -145 833 -111
rect 867 -145 901 -111
rect 935 -145 969 -111
rect 1003 -145 1037 -111
rect 1071 -145 1105 -111
rect 1139 -145 1173 -111
rect 1207 -145 1241 -111
rect 1275 -145 1309 -111
rect 1343 -145 1377 -111
rect 1411 -145 1445 -111
rect 1479 -145 1513 -111
rect 1547 -145 1581 -111
rect 1615 -145 1649 -111
rect 1683 -145 1717 -111
rect 1751 -145 1785 -111
rect 1819 -145 1853 -111
rect 1887 -145 1921 -111
rect 1955 -145 2000 -111
rect -2000 -161 2000 -145
<< polycont >>
rect -1955 -145 -1921 -111
rect -1887 -145 -1853 -111
rect -1819 -145 -1785 -111
rect -1751 -145 -1717 -111
rect -1683 -145 -1649 -111
rect -1615 -145 -1581 -111
rect -1547 -145 -1513 -111
rect -1479 -145 -1445 -111
rect -1411 -145 -1377 -111
rect -1343 -145 -1309 -111
rect -1275 -145 -1241 -111
rect -1207 -145 -1173 -111
rect -1139 -145 -1105 -111
rect -1071 -145 -1037 -111
rect -1003 -145 -969 -111
rect -935 -145 -901 -111
rect -867 -145 -833 -111
rect -799 -145 -765 -111
rect -731 -145 -697 -111
rect -663 -145 -629 -111
rect -595 -145 -561 -111
rect -527 -145 -493 -111
rect -459 -145 -425 -111
rect -391 -145 -357 -111
rect -323 -145 -289 -111
rect -255 -145 -221 -111
rect -187 -145 -153 -111
rect -119 -145 -85 -111
rect -51 -145 -17 -111
rect 17 -145 51 -111
rect 85 -145 119 -111
rect 153 -145 187 -111
rect 221 -145 255 -111
rect 289 -145 323 -111
rect 357 -145 391 -111
rect 425 -145 459 -111
rect 493 -145 527 -111
rect 561 -145 595 -111
rect 629 -145 663 -111
rect 697 -145 731 -111
rect 765 -145 799 -111
rect 833 -145 867 -111
rect 901 -145 935 -111
rect 969 -145 1003 -111
rect 1037 -145 1071 -111
rect 1105 -145 1139 -111
rect 1173 -145 1207 -111
rect 1241 -145 1275 -111
rect 1309 -145 1343 -111
rect 1377 -145 1411 -111
rect 1445 -145 1479 -111
rect 1513 -145 1547 -111
rect 1581 -145 1615 -111
rect 1649 -145 1683 -111
rect 1717 -145 1751 -111
rect 1785 -145 1819 -111
rect 1853 -145 1887 -111
rect 1921 -145 1955 -111
<< locali >>
rect -2160 214 -2057 248
rect -2023 214 -1989 248
rect -1955 214 -1921 248
rect -1887 214 -1853 248
rect -1819 214 -1785 248
rect -1751 214 -1717 248
rect -1683 214 -1649 248
rect -1615 214 -1581 248
rect -1547 214 -1513 248
rect -1479 214 -1445 248
rect -1411 214 -1377 248
rect -1343 214 -1309 248
rect -1275 214 -1241 248
rect -1207 214 -1173 248
rect -1139 214 -1105 248
rect -1071 214 -1037 248
rect -1003 214 -969 248
rect -935 214 -901 248
rect -867 214 -833 248
rect -799 214 -765 248
rect -731 214 -697 248
rect -663 214 -629 248
rect -595 214 -561 248
rect -527 214 -493 248
rect -459 214 -425 248
rect -391 214 -357 248
rect -323 214 -289 248
rect -255 214 -221 248
rect -187 214 -153 248
rect -119 214 -85 248
rect -51 214 -17 248
rect 17 214 51 248
rect 85 214 119 248
rect 153 214 187 248
rect 221 214 255 248
rect 289 214 323 248
rect 357 214 391 248
rect 425 214 459 248
rect 493 214 527 248
rect 561 214 595 248
rect 629 214 663 248
rect 697 214 731 248
rect 765 214 799 248
rect 833 214 867 248
rect 901 214 935 248
rect 969 214 1003 248
rect 1037 214 1071 248
rect 1105 214 1139 248
rect 1173 214 1207 248
rect 1241 214 1275 248
rect 1309 214 1343 248
rect 1377 214 1411 248
rect 1445 214 1479 248
rect 1513 214 1547 248
rect 1581 214 1615 248
rect 1649 214 1683 248
rect 1717 214 1751 248
rect 1785 214 1819 248
rect 1853 214 1887 248
rect 1921 214 1955 248
rect 1989 214 2023 248
rect 2057 214 2160 248
rect -2160 -214 -2126 214
rect -2046 121 -2012 140
rect -2046 53 -2012 55
rect -2046 17 -2012 19
rect -2046 -68 -2012 -49
rect 2012 121 2046 140
rect 2012 53 2046 55
rect 2012 17 2046 19
rect 2012 -68 2046 -49
rect -2000 -145 -1961 -111
rect -1921 -145 -1889 -111
rect -1853 -145 -1819 -111
rect -1783 -145 -1751 -111
rect -1711 -145 -1683 -111
rect -1639 -145 -1615 -111
rect -1567 -145 -1547 -111
rect -1495 -145 -1479 -111
rect -1423 -145 -1411 -111
rect -1351 -145 -1343 -111
rect -1279 -145 -1275 -111
rect -1173 -145 -1169 -111
rect -1105 -145 -1097 -111
rect -1037 -145 -1025 -111
rect -969 -145 -953 -111
rect -901 -145 -881 -111
rect -833 -145 -809 -111
rect -765 -145 -737 -111
rect -697 -145 -665 -111
rect -629 -145 -595 -111
rect -559 -145 -527 -111
rect -487 -145 -459 -111
rect -415 -145 -391 -111
rect -343 -145 -323 -111
rect -271 -145 -255 -111
rect -199 -145 -187 -111
rect -127 -145 -119 -111
rect -55 -145 -51 -111
rect 51 -145 55 -111
rect 119 -145 127 -111
rect 187 -145 199 -111
rect 255 -145 271 -111
rect 323 -145 343 -111
rect 391 -145 415 -111
rect 459 -145 487 -111
rect 527 -145 559 -111
rect 595 -145 629 -111
rect 665 -145 697 -111
rect 737 -145 765 -111
rect 809 -145 833 -111
rect 881 -145 901 -111
rect 953 -145 969 -111
rect 1025 -145 1037 -111
rect 1097 -145 1105 -111
rect 1169 -145 1173 -111
rect 1275 -145 1279 -111
rect 1343 -145 1351 -111
rect 1411 -145 1423 -111
rect 1479 -145 1495 -111
rect 1547 -145 1567 -111
rect 1615 -145 1639 -111
rect 1683 -145 1711 -111
rect 1751 -145 1783 -111
rect 1819 -145 1853 -111
rect 1889 -145 1921 -111
rect 1961 -145 2000 -111
rect 2126 -214 2160 214
rect -2160 -248 2160 -214
<< viali >>
rect -2046 87 -2012 89
rect -2046 55 -2012 87
rect -2046 -15 -2012 17
rect -2046 -17 -2012 -15
rect 2012 87 2046 89
rect 2012 55 2046 87
rect 2012 -15 2046 17
rect 2012 -17 2046 -15
rect -1961 -145 -1955 -111
rect -1955 -145 -1927 -111
rect -1889 -145 -1887 -111
rect -1887 -145 -1855 -111
rect -1817 -145 -1785 -111
rect -1785 -145 -1783 -111
rect -1745 -145 -1717 -111
rect -1717 -145 -1711 -111
rect -1673 -145 -1649 -111
rect -1649 -145 -1639 -111
rect -1601 -145 -1581 -111
rect -1581 -145 -1567 -111
rect -1529 -145 -1513 -111
rect -1513 -145 -1495 -111
rect -1457 -145 -1445 -111
rect -1445 -145 -1423 -111
rect -1385 -145 -1377 -111
rect -1377 -145 -1351 -111
rect -1313 -145 -1309 -111
rect -1309 -145 -1279 -111
rect -1241 -145 -1207 -111
rect -1169 -145 -1139 -111
rect -1139 -145 -1135 -111
rect -1097 -145 -1071 -111
rect -1071 -145 -1063 -111
rect -1025 -145 -1003 -111
rect -1003 -145 -991 -111
rect -953 -145 -935 -111
rect -935 -145 -919 -111
rect -881 -145 -867 -111
rect -867 -145 -847 -111
rect -809 -145 -799 -111
rect -799 -145 -775 -111
rect -737 -145 -731 -111
rect -731 -145 -703 -111
rect -665 -145 -663 -111
rect -663 -145 -631 -111
rect -593 -145 -561 -111
rect -561 -145 -559 -111
rect -521 -145 -493 -111
rect -493 -145 -487 -111
rect -449 -145 -425 -111
rect -425 -145 -415 -111
rect -377 -145 -357 -111
rect -357 -145 -343 -111
rect -305 -145 -289 -111
rect -289 -145 -271 -111
rect -233 -145 -221 -111
rect -221 -145 -199 -111
rect -161 -145 -153 -111
rect -153 -145 -127 -111
rect -89 -145 -85 -111
rect -85 -145 -55 -111
rect -17 -145 17 -111
rect 55 -145 85 -111
rect 85 -145 89 -111
rect 127 -145 153 -111
rect 153 -145 161 -111
rect 199 -145 221 -111
rect 221 -145 233 -111
rect 271 -145 289 -111
rect 289 -145 305 -111
rect 343 -145 357 -111
rect 357 -145 377 -111
rect 415 -145 425 -111
rect 425 -145 449 -111
rect 487 -145 493 -111
rect 493 -145 521 -111
rect 559 -145 561 -111
rect 561 -145 593 -111
rect 631 -145 663 -111
rect 663 -145 665 -111
rect 703 -145 731 -111
rect 731 -145 737 -111
rect 775 -145 799 -111
rect 799 -145 809 -111
rect 847 -145 867 -111
rect 867 -145 881 -111
rect 919 -145 935 -111
rect 935 -145 953 -111
rect 991 -145 1003 -111
rect 1003 -145 1025 -111
rect 1063 -145 1071 -111
rect 1071 -145 1097 -111
rect 1135 -145 1139 -111
rect 1139 -145 1169 -111
rect 1207 -145 1241 -111
rect 1279 -145 1309 -111
rect 1309 -145 1313 -111
rect 1351 -145 1377 -111
rect 1377 -145 1385 -111
rect 1423 -145 1445 -111
rect 1445 -145 1457 -111
rect 1495 -145 1513 -111
rect 1513 -145 1529 -111
rect 1567 -145 1581 -111
rect 1581 -145 1601 -111
rect 1639 -145 1649 -111
rect 1649 -145 1673 -111
rect 1711 -145 1717 -111
rect 1717 -145 1745 -111
rect 1783 -145 1785 -111
rect 1785 -145 1817 -111
rect 1855 -145 1887 -111
rect 1887 -145 1889 -111
rect 1927 -145 1955 -111
rect 1955 -145 1961 -111
<< metal1 >>
rect -2052 89 -2006 136
rect -2052 55 -2046 89
rect -2012 55 -2006 89
rect -2052 17 -2006 55
rect -2052 -17 -2046 17
rect -2012 -17 -2006 17
rect -2052 -64 -2006 -17
rect 2006 89 2052 136
rect 2006 55 2012 89
rect 2046 55 2052 89
rect 2006 17 2052 55
rect 2006 -17 2012 17
rect 2046 -17 2052 17
rect 2006 -64 2052 -17
rect -1996 -111 1996 -105
rect -1996 -145 -1961 -111
rect -1927 -145 -1889 -111
rect -1855 -145 -1817 -111
rect -1783 -145 -1745 -111
rect -1711 -145 -1673 -111
rect -1639 -145 -1601 -111
rect -1567 -145 -1529 -111
rect -1495 -145 -1457 -111
rect -1423 -145 -1385 -111
rect -1351 -145 -1313 -111
rect -1279 -145 -1241 -111
rect -1207 -145 -1169 -111
rect -1135 -145 -1097 -111
rect -1063 -145 -1025 -111
rect -991 -145 -953 -111
rect -919 -145 -881 -111
rect -847 -145 -809 -111
rect -775 -145 -737 -111
rect -703 -145 -665 -111
rect -631 -145 -593 -111
rect -559 -145 -521 -111
rect -487 -145 -449 -111
rect -415 -145 -377 -111
rect -343 -145 -305 -111
rect -271 -145 -233 -111
rect -199 -145 -161 -111
rect -127 -145 -89 -111
rect -55 -145 -17 -111
rect 17 -145 55 -111
rect 89 -145 127 -111
rect 161 -145 199 -111
rect 233 -145 271 -111
rect 305 -145 343 -111
rect 377 -145 415 -111
rect 449 -145 487 -111
rect 521 -145 559 -111
rect 593 -145 631 -111
rect 665 -145 703 -111
rect 737 -145 775 -111
rect 809 -145 847 -111
rect 881 -145 919 -111
rect 953 -145 991 -111
rect 1025 -145 1063 -111
rect 1097 -145 1135 -111
rect 1169 -145 1207 -111
rect 1241 -145 1279 -111
rect 1313 -145 1351 -111
rect 1385 -145 1423 -111
rect 1457 -145 1495 -111
rect 1529 -145 1567 -111
rect 1601 -145 1639 -111
rect 1673 -145 1711 -111
rect 1745 -145 1783 -111
rect 1817 -145 1855 -111
rect 1889 -145 1927 -111
rect 1961 -145 1996 -111
rect -1996 -151 1996 -145
<< properties >>
string FIXED_BBOX -2143 -231 2143 231
<< end >>
