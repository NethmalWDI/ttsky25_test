magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< error_s >>
rect -628 1740 -272 1868
rect -628 1700 -480 1740
rect -460 1700 -440 1740
rect -460 1620 -206 1700
rect -440 1584 -404 1620
<< nwell >>
rect -480 1700 4000 1740
rect -480 1620 -460 1700
rect -440 1620 4000 1700
rect -480 -1940 4000 1620
<< nsubdiff >>
rect -440 1677 3960 1700
rect -440 1643 -345 1677
rect -311 1643 -277 1677
rect -243 1643 -209 1677
rect -175 1643 -141 1677
rect -107 1643 -73 1677
rect -39 1643 -5 1677
rect 29 1643 63 1677
rect 97 1643 131 1677
rect 165 1643 199 1677
rect 233 1643 267 1677
rect 301 1643 335 1677
rect 369 1643 403 1677
rect 437 1643 471 1677
rect 505 1643 539 1677
rect 573 1643 607 1677
rect 641 1643 675 1677
rect 709 1643 743 1677
rect 777 1643 811 1677
rect 845 1643 879 1677
rect 913 1643 947 1677
rect 981 1643 1015 1677
rect 1049 1643 1083 1677
rect 1117 1643 1151 1677
rect 1185 1643 1219 1677
rect 1253 1643 1287 1677
rect 1321 1643 1355 1677
rect 1389 1643 1423 1677
rect 1457 1643 1491 1677
rect 1525 1643 1559 1677
rect 1593 1643 1627 1677
rect 1661 1643 1695 1677
rect 1729 1643 1763 1677
rect 1797 1643 1831 1677
rect 1865 1643 1899 1677
rect 1933 1643 1967 1677
rect 2001 1643 2035 1677
rect 2069 1643 2103 1677
rect 2137 1643 2171 1677
rect 2205 1643 2239 1677
rect 2273 1643 2307 1677
rect 2341 1643 2375 1677
rect 2409 1643 2443 1677
rect 2477 1643 2511 1677
rect 2545 1643 2579 1677
rect 2613 1643 2647 1677
rect 2681 1643 2715 1677
rect 2749 1643 2783 1677
rect 2817 1643 2851 1677
rect 2885 1643 2919 1677
rect 2953 1643 2987 1677
rect 3021 1643 3055 1677
rect 3089 1643 3123 1677
rect 3157 1643 3191 1677
rect 3225 1643 3259 1677
rect 3293 1643 3327 1677
rect 3361 1643 3395 1677
rect 3429 1643 3463 1677
rect 3497 1643 3531 1677
rect 3565 1643 3599 1677
rect 3633 1643 3667 1677
rect 3701 1643 3735 1677
rect 3769 1643 3803 1677
rect 3837 1643 3871 1677
rect 3905 1643 3960 1677
rect -440 1620 3960 1643
rect -440 -1860 -400 1620
rect 3920 -1860 3960 1620
rect -440 -1900 3960 -1860
<< nsubdiffcont >>
rect -345 1643 -311 1677
rect -277 1643 -243 1677
rect -209 1643 -175 1677
rect -141 1643 -107 1677
rect -73 1643 -39 1677
rect -5 1643 29 1677
rect 63 1643 97 1677
rect 131 1643 165 1677
rect 199 1643 233 1677
rect 267 1643 301 1677
rect 335 1643 369 1677
rect 403 1643 437 1677
rect 471 1643 505 1677
rect 539 1643 573 1677
rect 607 1643 641 1677
rect 675 1643 709 1677
rect 743 1643 777 1677
rect 811 1643 845 1677
rect 879 1643 913 1677
rect 947 1643 981 1677
rect 1015 1643 1049 1677
rect 1083 1643 1117 1677
rect 1151 1643 1185 1677
rect 1219 1643 1253 1677
rect 1287 1643 1321 1677
rect 1355 1643 1389 1677
rect 1423 1643 1457 1677
rect 1491 1643 1525 1677
rect 1559 1643 1593 1677
rect 1627 1643 1661 1677
rect 1695 1643 1729 1677
rect 1763 1643 1797 1677
rect 1831 1643 1865 1677
rect 1899 1643 1933 1677
rect 1967 1643 2001 1677
rect 2035 1643 2069 1677
rect 2103 1643 2137 1677
rect 2171 1643 2205 1677
rect 2239 1643 2273 1677
rect 2307 1643 2341 1677
rect 2375 1643 2409 1677
rect 2443 1643 2477 1677
rect 2511 1643 2545 1677
rect 2579 1643 2613 1677
rect 2647 1643 2681 1677
rect 2715 1643 2749 1677
rect 2783 1643 2817 1677
rect 2851 1643 2885 1677
rect 2919 1643 2953 1677
rect 2987 1643 3021 1677
rect 3055 1643 3089 1677
rect 3123 1643 3157 1677
rect 3191 1643 3225 1677
rect 3259 1643 3293 1677
rect 3327 1643 3361 1677
rect 3395 1643 3429 1677
rect 3463 1643 3497 1677
rect 3531 1643 3565 1677
rect 3599 1643 3633 1677
rect 3667 1643 3701 1677
rect 3735 1643 3769 1677
rect 3803 1643 3837 1677
rect 3871 1643 3905 1677
<< locali >>
rect -440 1677 3960 1700
rect -440 1643 -345 1677
rect -291 1643 -277 1677
rect -219 1643 -209 1677
rect -147 1643 -141 1677
rect -75 1643 -73 1677
rect -39 1643 -37 1677
rect 29 1643 35 1677
rect 97 1643 107 1677
rect 165 1643 179 1677
rect 233 1643 251 1677
rect 301 1643 323 1677
rect 369 1643 395 1677
rect 437 1643 467 1677
rect 505 1643 539 1677
rect 573 1643 607 1677
rect 645 1643 675 1677
rect 717 1643 743 1677
rect 789 1643 811 1677
rect 861 1643 879 1677
rect 933 1643 947 1677
rect 1005 1643 1015 1677
rect 1077 1643 1083 1677
rect 1149 1643 1151 1677
rect 1185 1643 1187 1677
rect 1253 1643 1259 1677
rect 1321 1643 1331 1677
rect 1389 1643 1403 1677
rect 1457 1643 1475 1677
rect 1525 1643 1547 1677
rect 1593 1643 1619 1677
rect 1661 1643 1691 1677
rect 1729 1643 1763 1677
rect 1797 1643 1831 1677
rect 1869 1643 1899 1677
rect 1941 1643 1967 1677
rect 2013 1643 2035 1677
rect 2085 1643 2103 1677
rect 2157 1643 2171 1677
rect 2229 1643 2239 1677
rect 2301 1643 2307 1677
rect 2373 1643 2375 1677
rect 2409 1643 2411 1677
rect 2477 1643 2483 1677
rect 2545 1643 2555 1677
rect 2613 1643 2627 1677
rect 2681 1643 2699 1677
rect 2749 1643 2771 1677
rect 2817 1643 2843 1677
rect 2885 1643 2915 1677
rect 2953 1643 2987 1677
rect 3021 1643 3055 1677
rect 3093 1643 3123 1677
rect 3165 1643 3191 1677
rect 3237 1643 3259 1677
rect 3309 1643 3327 1677
rect 3381 1643 3395 1677
rect 3453 1643 3463 1677
rect 3525 1643 3531 1677
rect 3597 1643 3599 1677
rect 3633 1643 3635 1677
rect 3701 1643 3707 1677
rect 3769 1643 3779 1677
rect 3837 1643 3851 1677
rect 3905 1643 3960 1677
rect -440 1620 3960 1643
rect -440 -1860 -400 1620
rect 3920 -1860 3960 1620
rect -440 -1900 3960 -1860
<< viali >>
rect -325 1643 -311 1677
rect -311 1643 -291 1677
rect -253 1643 -243 1677
rect -243 1643 -219 1677
rect -181 1643 -175 1677
rect -175 1643 -147 1677
rect -109 1643 -107 1677
rect -107 1643 -75 1677
rect -37 1643 -5 1677
rect -5 1643 -3 1677
rect 35 1643 63 1677
rect 63 1643 69 1677
rect 107 1643 131 1677
rect 131 1643 141 1677
rect 179 1643 199 1677
rect 199 1643 213 1677
rect 251 1643 267 1677
rect 267 1643 285 1677
rect 323 1643 335 1677
rect 335 1643 357 1677
rect 395 1643 403 1677
rect 403 1643 429 1677
rect 467 1643 471 1677
rect 471 1643 501 1677
rect 539 1643 573 1677
rect 611 1643 641 1677
rect 641 1643 645 1677
rect 683 1643 709 1677
rect 709 1643 717 1677
rect 755 1643 777 1677
rect 777 1643 789 1677
rect 827 1643 845 1677
rect 845 1643 861 1677
rect 899 1643 913 1677
rect 913 1643 933 1677
rect 971 1643 981 1677
rect 981 1643 1005 1677
rect 1043 1643 1049 1677
rect 1049 1643 1077 1677
rect 1115 1643 1117 1677
rect 1117 1643 1149 1677
rect 1187 1643 1219 1677
rect 1219 1643 1221 1677
rect 1259 1643 1287 1677
rect 1287 1643 1293 1677
rect 1331 1643 1355 1677
rect 1355 1643 1365 1677
rect 1403 1643 1423 1677
rect 1423 1643 1437 1677
rect 1475 1643 1491 1677
rect 1491 1643 1509 1677
rect 1547 1643 1559 1677
rect 1559 1643 1581 1677
rect 1619 1643 1627 1677
rect 1627 1643 1653 1677
rect 1691 1643 1695 1677
rect 1695 1643 1725 1677
rect 1763 1643 1797 1677
rect 1835 1643 1865 1677
rect 1865 1643 1869 1677
rect 1907 1643 1933 1677
rect 1933 1643 1941 1677
rect 1979 1643 2001 1677
rect 2001 1643 2013 1677
rect 2051 1643 2069 1677
rect 2069 1643 2085 1677
rect 2123 1643 2137 1677
rect 2137 1643 2157 1677
rect 2195 1643 2205 1677
rect 2205 1643 2229 1677
rect 2267 1643 2273 1677
rect 2273 1643 2301 1677
rect 2339 1643 2341 1677
rect 2341 1643 2373 1677
rect 2411 1643 2443 1677
rect 2443 1643 2445 1677
rect 2483 1643 2511 1677
rect 2511 1643 2517 1677
rect 2555 1643 2579 1677
rect 2579 1643 2589 1677
rect 2627 1643 2647 1677
rect 2647 1643 2661 1677
rect 2699 1643 2715 1677
rect 2715 1643 2733 1677
rect 2771 1643 2783 1677
rect 2783 1643 2805 1677
rect 2843 1643 2851 1677
rect 2851 1643 2877 1677
rect 2915 1643 2919 1677
rect 2919 1643 2949 1677
rect 2987 1643 3021 1677
rect 3059 1643 3089 1677
rect 3089 1643 3093 1677
rect 3131 1643 3157 1677
rect 3157 1643 3165 1677
rect 3203 1643 3225 1677
rect 3225 1643 3237 1677
rect 3275 1643 3293 1677
rect 3293 1643 3309 1677
rect 3347 1643 3361 1677
rect 3361 1643 3381 1677
rect 3419 1643 3429 1677
rect 3429 1643 3453 1677
rect 3491 1643 3497 1677
rect 3497 1643 3525 1677
rect 3563 1643 3565 1677
rect 3565 1643 3597 1677
rect 3635 1643 3667 1677
rect 3667 1643 3669 1677
rect 3707 1643 3735 1677
rect 3735 1643 3741 1677
rect 3779 1643 3803 1677
rect 3803 1643 3813 1677
rect 3851 1643 3871 1677
rect 3871 1643 3885 1677
<< metal1 >>
rect -440 1677 3960 1700
rect -440 1643 -325 1677
rect -291 1643 -253 1677
rect -219 1643 -181 1677
rect -147 1643 -109 1677
rect -75 1643 -37 1677
rect -3 1643 35 1677
rect 69 1643 107 1677
rect 141 1643 179 1677
rect 213 1643 251 1677
rect 285 1643 323 1677
rect 357 1643 395 1677
rect 429 1643 467 1677
rect 501 1643 539 1677
rect 573 1643 611 1677
rect 645 1643 683 1677
rect 717 1643 755 1677
rect 789 1643 827 1677
rect 861 1643 899 1677
rect 933 1643 971 1677
rect 1005 1643 1043 1677
rect 1077 1643 1115 1677
rect 1149 1643 1187 1677
rect 1221 1643 1259 1677
rect 1293 1643 1331 1677
rect 1365 1643 1403 1677
rect 1437 1643 1475 1677
rect 1509 1643 1547 1677
rect 1581 1643 1619 1677
rect 1653 1643 1691 1677
rect 1725 1643 1763 1677
rect 1797 1643 1835 1677
rect 1869 1643 1907 1677
rect 1941 1643 1979 1677
rect 2013 1643 2051 1677
rect 2085 1643 2123 1677
rect 2157 1643 2195 1677
rect 2229 1643 2267 1677
rect 2301 1643 2339 1677
rect 2373 1643 2411 1677
rect 2445 1643 2483 1677
rect 2517 1643 2555 1677
rect 2589 1643 2627 1677
rect 2661 1643 2699 1677
rect 2733 1643 2771 1677
rect 2805 1643 2843 1677
rect 2877 1643 2915 1677
rect 2949 1643 2987 1677
rect 3021 1643 3059 1677
rect 3093 1643 3131 1677
rect 3165 1643 3203 1677
rect 3237 1643 3275 1677
rect 3309 1643 3347 1677
rect 3381 1643 3419 1677
rect 3453 1643 3491 1677
rect 3525 1643 3563 1677
rect 3597 1643 3635 1677
rect 3669 1643 3707 1677
rect 3741 1643 3779 1677
rect 3813 1643 3851 1677
rect 3885 1643 3960 1677
rect -440 1620 3960 1643
rect 0 1500 3860 1620
rect 0 1180 60 1500
rect 300 1260 360 1500
rect -150 1156 -70 1160
rect -150 1104 -136 1156
rect -84 1104 -70 1156
rect -150 1100 -70 1104
rect 0 1100 380 1180
rect -390 -4 -310 0
rect -390 -56 -376 -4
rect -324 -56 -310 -4
rect -390 -60 -310 -56
rect -380 -70 -320 -60
rect -270 -124 -190 -120
rect -270 -176 -256 -124
rect -204 -176 -190 -124
rect -270 -180 -190 -176
rect -260 -190 -200 -180
rect -140 -240 -80 1100
rect 0 960 60 1100
rect 0 400 80 960
rect 0 -240 60 400
rect 300 60 380 1100
rect -150 -244 -70 -240
rect -150 -296 -136 -244
rect -84 -296 -70 -244
rect -150 -300 -70 -296
rect 0 -300 360 -240
rect -140 -310 -80 -300
rect 0 -1440 60 -300
rect 300 -1320 360 -300
rect 500 -1320 560 1500
rect 800 1260 860 1500
rect 620 1166 760 1170
rect 620 1114 632 1166
rect 684 1114 696 1166
rect 748 1114 760 1166
rect 620 1110 760 1114
rect 800 -120 860 1040
rect 790 -124 870 -120
rect 790 -176 804 -124
rect 856 -176 870 -124
rect 790 -180 870 -176
rect 620 -234 760 -230
rect 620 -286 632 -234
rect 684 -286 696 -234
rect 748 -286 760 -234
rect 620 -290 760 -286
rect 820 -762 940 -740
rect 820 -814 864 -762
rect 916 -814 940 -762
rect 820 -826 940 -814
rect 820 -878 864 -826
rect 916 -878 940 -826
rect 820 -900 940 -878
rect 1000 -1320 1060 1500
rect 1300 1260 1360 1500
rect 1120 1166 1260 1170
rect 1120 1114 1132 1166
rect 1184 1114 1196 1166
rect 1248 1114 1260 1166
rect 1120 1110 1260 1114
rect 1300 0 1360 1060
rect 1290 -4 1370 0
rect 1290 -56 1304 -4
rect 1356 -56 1370 -4
rect 1290 -60 1370 -56
rect 1120 -234 1260 -230
rect 1120 -286 1132 -234
rect 1184 -286 1196 -234
rect 1248 -286 1260 -234
rect 1120 -290 1260 -286
rect 1500 -240 1560 1500
rect 1800 1260 1860 1500
rect 1620 1166 1760 1170
rect 1620 1114 1632 1166
rect 1684 1114 1696 1166
rect 1748 1160 1760 1166
rect 2000 1160 2060 1500
rect 2300 1260 2360 1500
rect 1748 1114 1860 1160
rect 1620 1110 1860 1114
rect 1660 1100 1860 1110
rect 1800 640 1860 1100
rect 2000 1100 2360 1160
rect 1800 618 1940 640
rect 1800 566 1864 618
rect 1916 566 1940 618
rect 1800 554 1940 566
rect 1800 502 1864 554
rect 1916 502 1940 554
rect 1800 480 1940 502
rect 1500 -300 1860 -240
rect 1320 -762 1440 -740
rect 1320 -814 1364 -762
rect 1416 -814 1440 -762
rect 1320 -826 1440 -814
rect 1320 -878 1364 -826
rect 1416 -878 1440 -826
rect 1320 -900 1440 -878
rect 1500 -1320 1560 -300
rect 1800 -1340 1860 -300
rect 2000 -1320 2060 1100
rect 2300 60 2360 1100
rect 2120 -234 2260 -230
rect 2120 -286 2132 -234
rect 2184 -286 2196 -234
rect 2248 -240 2260 -234
rect 2248 -286 2360 -240
rect 2120 -290 2360 -286
rect 2140 -300 2360 -290
rect 2300 -760 2360 -300
rect 2300 -780 2440 -760
rect 2320 -782 2440 -780
rect 2320 -834 2364 -782
rect 2416 -834 2440 -782
rect 2320 -846 2440 -834
rect 2320 -898 2364 -846
rect 2416 -898 2440 -846
rect 2320 -920 2440 -898
rect 2500 -1320 2560 1500
rect 2800 1260 2860 1500
rect 2620 1166 2760 1170
rect 2620 1114 2632 1166
rect 2684 1114 2696 1166
rect 2748 1114 2760 1166
rect 2620 1110 2760 1114
rect 2820 618 2940 640
rect 2820 566 2864 618
rect 2916 566 2940 618
rect 2820 554 2940 566
rect 2820 502 2864 554
rect 2916 502 2940 554
rect 2820 480 2940 502
rect 2810 -4 2890 0
rect 2810 -56 2824 -4
rect 2876 -56 2890 -4
rect 2810 -60 2890 -56
rect 2620 -234 2760 -230
rect 2620 -286 2632 -234
rect 2684 -286 2696 -234
rect 2748 -286 2760 -234
rect 2620 -290 2760 -286
rect 2820 -1340 2880 -60
rect 3000 -1320 3060 1500
rect 3300 1260 3360 1500
rect 3120 1166 3260 1170
rect 3120 1114 3132 1166
rect 3184 1114 3196 1166
rect 3248 1114 3260 1166
rect 3120 1110 3260 1114
rect 3500 1160 3560 1500
rect 3800 1260 3860 1500
rect 3500 1100 3860 1160
rect 3320 618 3440 640
rect 3320 566 3364 618
rect 3416 566 3440 618
rect 3320 554 3440 566
rect 3320 502 3364 554
rect 3416 502 3440 554
rect 3320 480 3440 502
rect 3310 -124 3390 -120
rect 3310 -176 3324 -124
rect 3376 -176 3390 -124
rect 3310 -180 3390 -176
rect 3120 -234 3260 -230
rect 3120 -286 3132 -234
rect 3184 -286 3196 -234
rect 3248 -286 3260 -234
rect 3120 -290 3260 -286
rect 3320 -1340 3380 -180
rect 3500 -240 3560 1100
rect 3800 60 3860 1100
rect 3500 -300 3860 -240
rect 3500 -1300 3560 -300
rect 3800 -1340 3860 -300
rect 0 -1500 3860 -1440
rect 0 -1740 60 -1500
rect 300 -1740 360 -1500
rect 520 -1740 580 -1500
rect 800 -1740 860 -1500
rect 1040 -1740 1100 -1500
rect 1320 -1740 1380 -1500
rect 1540 -1740 1600 -1500
rect 1800 -1740 1860 -1500
rect 2020 -1740 2080 -1500
rect 2300 -1740 2360 -1500
rect 2540 -1740 2600 -1500
rect 2800 -1740 2860 -1500
rect 3020 -1740 3080 -1500
rect 3300 -1740 3360 -1500
rect 3520 -1740 3580 -1500
rect 3800 -1740 3860 -1500
<< via1 >>
rect -136 1104 -84 1156
rect -376 -56 -324 -4
rect -256 -176 -204 -124
rect -136 -296 -84 -244
rect 632 1114 684 1166
rect 696 1114 748 1166
rect 804 -176 856 -124
rect 632 -286 684 -234
rect 696 -286 748 -234
rect 864 -814 916 -762
rect 864 -878 916 -826
rect 1132 1114 1184 1166
rect 1196 1114 1248 1166
rect 1304 -56 1356 -4
rect 1132 -286 1184 -234
rect 1196 -286 1248 -234
rect 1632 1114 1684 1166
rect 1696 1114 1748 1166
rect 1864 566 1916 618
rect 1864 502 1916 554
rect 1364 -814 1416 -762
rect 1364 -878 1416 -826
rect 2132 -286 2184 -234
rect 2196 -286 2248 -234
rect 2364 -834 2416 -782
rect 2364 -898 2416 -846
rect 2632 1114 2684 1166
rect 2696 1114 2748 1166
rect 2864 566 2916 618
rect 2864 502 2916 554
rect 2824 -56 2876 -4
rect 2632 -286 2684 -234
rect 2696 -286 2748 -234
rect 3132 1114 3184 1166
rect 3196 1114 3248 1166
rect 3364 566 3416 618
rect 3364 502 3416 554
rect 3324 -176 3376 -124
rect 3132 -286 3184 -234
rect 3196 -286 3248 -234
<< metal2 >>
rect -140 1160 -80 1170
rect 630 1166 750 1180
rect 630 1160 632 1166
rect -140 1156 632 1160
rect -140 1104 -136 1156
rect -84 1114 632 1156
rect 684 1114 696 1166
rect 748 1160 750 1166
rect 1130 1166 1250 1180
rect 1130 1160 1132 1166
rect 748 1114 1132 1160
rect 1184 1114 1196 1166
rect 1248 1160 1250 1166
rect 1630 1166 1750 1180
rect 1630 1160 1632 1166
rect 1248 1114 1632 1160
rect 1684 1114 1696 1166
rect 1748 1160 1750 1166
rect 2630 1166 2750 1180
rect 2630 1160 2632 1166
rect 1748 1114 2632 1160
rect 2684 1114 2696 1166
rect 2748 1160 2750 1166
rect 3130 1166 3250 1180
rect 3130 1160 3132 1166
rect 2748 1114 3132 1160
rect 3184 1114 3196 1166
rect 3248 1160 3250 1166
rect 3248 1114 3940 1160
rect -84 1104 3940 1114
rect -140 1100 3940 1104
rect -140 1090 -80 1100
rect 1860 618 1920 630
rect 1860 588 1864 618
rect 1916 588 1920 618
rect 1860 532 1862 588
rect 1918 532 1920 588
rect 1860 502 1864 532
rect 1916 502 1920 532
rect 1860 490 1920 502
rect 2860 618 2920 630
rect 2860 588 2864 618
rect 2916 588 2920 618
rect 2860 532 2862 588
rect 2918 532 2920 588
rect 2860 502 2864 532
rect 2916 502 2920 532
rect 2860 490 2920 502
rect 3360 618 3420 630
rect 3360 588 3364 618
rect 3416 588 3420 618
rect 3360 532 3362 588
rect 3418 532 3420 588
rect 3360 502 3364 532
rect 3416 502 3420 532
rect 3360 490 3420 502
rect -380 0 -320 10
rect 1300 0 1360 10
rect 2820 0 2880 10
rect -450 -4 2880 0
rect -450 -12 -376 -4
rect -450 -68 -438 -12
rect -382 -56 -376 -12
rect -324 -56 1304 -4
rect 1356 -56 2824 -4
rect 2876 -56 2880 -4
rect -382 -60 2880 -56
rect -382 -68 -320 -60
rect -450 -70 -320 -68
rect 1300 -70 1360 -60
rect 2820 -70 2880 -60
rect -450 -80 -370 -70
rect -260 -120 -200 -110
rect 800 -120 860 -110
rect 3320 -120 3380 -110
rect -310 -124 3380 -120
rect -310 -132 -256 -124
rect -310 -188 -298 -132
rect -204 -176 804 -124
rect 856 -176 3324 -124
rect 3376 -176 3380 -124
rect -242 -180 3380 -176
rect -242 -188 -200 -180
rect -310 -190 -200 -188
rect 800 -190 860 -180
rect 3320 -190 3380 -180
rect -310 -200 -230 -190
rect -140 -240 -80 -230
rect 630 -234 750 -220
rect 630 -240 632 -234
rect -170 -244 632 -240
rect -170 -252 -136 -244
rect -170 -308 -158 -252
rect -84 -286 632 -244
rect 684 -286 696 -234
rect 748 -240 750 -234
rect 1130 -234 1250 -220
rect 1130 -240 1132 -234
rect 748 -286 1132 -240
rect 1184 -286 1196 -234
rect 1248 -240 1250 -234
rect 2130 -234 2250 -220
rect 2130 -240 2132 -234
rect 1248 -286 2132 -240
rect 2184 -286 2196 -234
rect 2248 -240 2250 -234
rect 2630 -234 2750 -220
rect 2630 -240 2632 -234
rect 2248 -286 2632 -240
rect 2684 -286 2696 -234
rect 2748 -240 2750 -234
rect 3130 -234 3250 -220
rect 3130 -240 3132 -234
rect 2748 -286 3132 -240
rect 3184 -286 3196 -234
rect 3248 -240 3250 -234
rect 3248 -286 3920 -240
rect -84 -296 3920 -286
rect -102 -300 3920 -296
rect -102 -308 -80 -300
rect -170 -310 -80 -308
rect -170 -320 -90 -310
rect 860 -762 920 -750
rect 860 -792 864 -762
rect 916 -792 920 -762
rect 860 -848 862 -792
rect 918 -848 920 -792
rect 860 -878 864 -848
rect 916 -878 920 -848
rect 860 -890 920 -878
rect 1360 -762 1420 -750
rect 1360 -792 1364 -762
rect 1416 -792 1420 -762
rect 1360 -848 1362 -792
rect 1418 -848 1420 -792
rect 1360 -878 1364 -848
rect 1416 -878 1420 -848
rect 1360 -890 1420 -878
rect 2360 -782 2420 -770
rect 2360 -812 2364 -782
rect 2416 -812 2420 -782
rect 2360 -868 2362 -812
rect 2418 -868 2420 -812
rect 2360 -898 2364 -868
rect 2416 -898 2420 -868
rect 2360 -910 2420 -898
rect 1860 -1800 1940 -1790
rect 2360 -1800 2440 -1790
rect 1860 -1802 2440 -1800
rect 1860 -1858 1872 -1802
rect 1928 -1858 2372 -1802
rect 2428 -1858 2440 -1802
rect 1860 -1860 2440 -1858
rect 1860 -1870 1940 -1860
rect 2360 -1870 2440 -1860
rect -30 -1922 2950 -1910
rect -30 -1978 -18 -1922
rect 38 -1978 1372 -1922
rect 1428 -1978 2872 -1922
rect 2928 -1978 2950 -1922
rect -30 -1990 2950 -1978
rect 110 -2042 3450 -2030
rect 110 -2098 122 -2042
rect 178 -2098 872 -2042
rect 928 -2098 3372 -2042
rect 3428 -2098 3450 -2042
rect 110 -2110 3450 -2098
<< via2 >>
rect 1862 566 1864 588
rect 1864 566 1916 588
rect 1916 566 1918 588
rect 1862 554 1918 566
rect 1862 532 1864 554
rect 1864 532 1916 554
rect 1916 532 1918 554
rect 2862 566 2864 588
rect 2864 566 2916 588
rect 2916 566 2918 588
rect 2862 554 2918 566
rect 2862 532 2864 554
rect 2864 532 2916 554
rect 2916 532 2918 554
rect 3362 566 3364 588
rect 3364 566 3416 588
rect 3416 566 3418 588
rect 3362 554 3418 566
rect 3362 532 3364 554
rect 3364 532 3416 554
rect 3416 532 3418 554
rect -438 -68 -382 -12
rect -298 -176 -256 -132
rect -256 -176 -242 -132
rect -298 -188 -242 -176
rect -158 -296 -136 -252
rect -136 -296 -102 -252
rect -158 -308 -102 -296
rect 862 -814 864 -792
rect 864 -814 916 -792
rect 916 -814 918 -792
rect 862 -826 918 -814
rect 862 -848 864 -826
rect 864 -848 916 -826
rect 916 -848 918 -826
rect 1362 -814 1364 -792
rect 1364 -814 1416 -792
rect 1416 -814 1418 -792
rect 1362 -826 1418 -814
rect 1362 -848 1364 -826
rect 1364 -848 1416 -826
rect 1416 -848 1418 -826
rect 2362 -834 2364 -812
rect 2364 -834 2416 -812
rect 2416 -834 2418 -812
rect 2362 -846 2418 -834
rect 2362 -868 2364 -846
rect 2364 -868 2416 -846
rect 2416 -868 2418 -846
rect 1872 -1858 1928 -1802
rect 2372 -1858 2428 -1802
rect -18 -1978 38 -1922
rect 1372 -1978 1428 -1922
rect 2872 -1978 2928 -1922
rect 122 -2098 178 -2042
rect 872 -2098 928 -2042
rect 3372 -2098 3428 -2042
<< metal3 >>
rect 1860 625 1940 640
rect 2860 625 2940 640
rect 3360 625 3440 640
rect 1850 588 1940 625
rect 1850 532 1862 588
rect 1918 532 1940 588
rect 1850 495 1940 532
rect 2850 588 2940 625
rect 2850 532 2862 588
rect 2918 532 2940 588
rect 2850 495 2940 532
rect 3350 588 3440 625
rect 3350 532 3362 588
rect 3418 532 3440 588
rect 3350 495 3440 532
rect -450 -12 -370 0
rect -450 -68 -438 -12
rect -382 -68 -370 -12
rect -450 -2090 -370 -68
rect -310 -132 -230 -120
rect -310 -188 -298 -132
rect -242 -188 -230 -132
rect -310 -2130 -230 -188
rect -170 -252 -90 -240
rect -170 -308 -158 -252
rect -102 -308 -90 -252
rect -170 -2110 -90 -308
rect 860 -755 940 -740
rect 1360 -755 1440 -740
rect 850 -792 940 -755
rect 850 -848 862 -792
rect 918 -848 940 -792
rect 850 -885 940 -848
rect 1350 -792 1440 -755
rect 1350 -848 1362 -792
rect 1418 -848 1440 -792
rect 1350 -885 1440 -848
rect -30 -1922 50 -1910
rect -30 -1978 -18 -1922
rect 38 -1978 50 -1922
rect -30 -2120 50 -1978
rect 110 -2042 190 -2030
rect 860 -2035 940 -885
rect 1360 -1915 1440 -885
rect 1860 -1795 1940 495
rect 2360 -775 2440 -760
rect 2350 -812 2440 -775
rect 2350 -868 2362 -812
rect 2418 -868 2440 -812
rect 2350 -905 2440 -868
rect 2360 -1340 2440 -905
rect 2300 -1795 2440 -1340
rect 1850 -1802 1950 -1795
rect 2300 -1800 2450 -1795
rect 1850 -1858 1872 -1802
rect 1928 -1858 1950 -1802
rect 1850 -1865 1950 -1858
rect 2350 -1802 2450 -1800
rect 2350 -1858 2372 -1802
rect 2428 -1858 2450 -1802
rect 2350 -1865 2450 -1858
rect 2860 -1915 2940 495
rect 1350 -1922 1450 -1915
rect 1350 -1978 1372 -1922
rect 1428 -1978 1450 -1922
rect 1350 -1985 1450 -1978
rect 2850 -1922 2950 -1915
rect 2850 -1978 2872 -1922
rect 2928 -1978 2950 -1922
rect 2850 -1985 2950 -1978
rect 3360 -2035 3440 495
rect 110 -2098 122 -2042
rect 178 -2098 190 -2042
rect 110 -2220 190 -2098
rect 850 -2042 950 -2035
rect 850 -2098 872 -2042
rect 928 -2098 950 -2042
rect 850 -2105 950 -2098
rect 3350 -2042 3450 -2035
rect 3350 -2098 3372 -2042
rect 3428 -2098 3450 -2042
rect 3350 -2105 3450 -2098
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_0
timestamp 1757161594
transform 1 0 2194 0 1 -1602
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_1
timestamp 1757161594
transform 1 0 194 0 1 1398
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_2
timestamp 1757161594
transform 1 0 3194 0 1 -1602
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_3
timestamp 1757161594
transform 1 0 2694 0 1 -1602
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_4
timestamp 1757161594
transform 1 0 194 0 1 -1602
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_5
timestamp 1757161594
transform 1 0 1694 0 1 -1602
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_6
timestamp 1757161594
transform 1 0 1194 0 1 -1602
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_7
timestamp 1757161594
transform 1 0 694 0 1 -1602
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_8
timestamp 1757161594
transform 1 0 3694 0 1 -1602
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_9
timestamp 1757161594
transform 1 0 3694 0 1 1398
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_10
timestamp 1757161594
transform 1 0 3194 0 1 1398
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_11
timestamp 1757161594
transform 1 0 2694 0 1 1398
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_12
timestamp 1757161594
transform 1 0 2194 0 1 1398
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_13
timestamp 1757161594
transform 1 0 1694 0 1 1398
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_14
timestamp 1757161594
transform 1 0 1194 0 1 1398
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_J8833D  sky130_fd_pr__pfet_01v8_lvt_J8833D_15
timestamp 1757161594
transform 1 0 694 0 1 1398
box -194 -198 194 164
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_0
timestamp 1757161594
transform 1 0 1194 0 1 -802
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_1
timestamp 1757161594
transform 1 0 194 0 1 598
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_2
timestamp 1757161594
transform 1 0 694 0 1 598
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_3
timestamp 1757161594
transform 1 0 1194 0 1 598
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_4
timestamp 1757161594
transform 1 0 1694 0 1 598
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_5
timestamp 1757161594
transform 1 0 2194 0 1 598
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_6
timestamp 1757161594
transform 1 0 2694 0 1 598
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_7
timestamp 1757161594
transform 1 0 3194 0 1 598
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_8
timestamp 1757161594
transform 1 0 3694 0 1 598
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_9
timestamp 1757161594
transform 1 0 194 0 1 -802
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_10
timestamp 1757161594
transform 1 0 694 0 1 -802
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_11
timestamp 1757161594
transform 1 0 2694 0 1 -802
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_12
timestamp 1757161594
transform 1 0 1694 0 1 -802
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_13
timestamp 1757161594
transform 1 0 2194 0 1 -802
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_14
timestamp 1757161594
transform 1 0 3694 0 1 -802
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_U8838H  sky130_fd_pr__pfet_01v8_lvt_U8838H_15
timestamp 1757161594
transform 1 0 3194 0 1 -802
box -194 -598 194 564
<< end >>
