magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< error_s >>
rect 6040 -2382 6120 -2370
rect 6040 -2438 6052 -2382
rect 6040 -2450 6120 -2438
<< pwell >>
rect -583 2967 5933 3053
rect -583 -2434 -497 2967
rect 5847 2636 5933 2967
rect 5544 2394 5933 2636
rect -583 -2837 -234 -2434
rect 5847 -2837 5933 2394
rect -583 -2923 5933 -2837
<< psubdiff >>
rect -557 2993 -470 3027
rect -436 2993 -402 3027
rect -368 2993 -334 3027
rect -300 2993 -266 3027
rect -232 2993 -198 3027
rect -164 2993 -130 3027
rect -96 2993 -62 3027
rect -28 2993 6 3027
rect 40 2993 74 3027
rect 108 2993 142 3027
rect 176 2993 210 3027
rect 244 2993 278 3027
rect 312 2993 346 3027
rect 380 2993 414 3027
rect 448 2993 482 3027
rect 516 2993 550 3027
rect 584 2993 618 3027
rect 652 2993 686 3027
rect 720 2993 754 3027
rect 788 2993 822 3027
rect 856 2993 890 3027
rect 924 2993 958 3027
rect 992 2993 1026 3027
rect 1060 2993 1094 3027
rect 1128 2993 1162 3027
rect 1196 2993 1230 3027
rect 1264 2993 1298 3027
rect 1332 2993 1366 3027
rect 1400 2993 1434 3027
rect 1468 2993 1502 3027
rect 1536 2993 1570 3027
rect 1604 2993 1638 3027
rect 1672 2993 1706 3027
rect 1740 2993 1774 3027
rect 1808 2993 1842 3027
rect 1876 2993 1910 3027
rect 1944 2993 1978 3027
rect 2012 2993 2046 3027
rect 2080 2993 2114 3027
rect 2148 2993 2182 3027
rect 2216 2993 2250 3027
rect 2284 2993 2318 3027
rect 2352 2993 2386 3027
rect 2420 2993 2454 3027
rect 2488 2993 2522 3027
rect 2556 2993 2590 3027
rect 2624 2993 2658 3027
rect 2692 2993 2726 3027
rect 2760 2993 2794 3027
rect 2828 2993 2862 3027
rect 2896 2993 2930 3027
rect 2964 2993 2998 3027
rect 3032 2993 3066 3027
rect 3100 2993 3134 3027
rect 3168 2993 3202 3027
rect 3236 2993 3270 3027
rect 3304 2993 3338 3027
rect 3372 2993 3406 3027
rect 3440 2993 3474 3027
rect 3508 2993 3542 3027
rect 3576 2993 3610 3027
rect 3644 2993 3678 3027
rect 3712 2993 3746 3027
rect 3780 2993 3814 3027
rect 3848 2993 3882 3027
rect 3916 2993 3950 3027
rect 3984 2993 4018 3027
rect 4052 2993 4086 3027
rect 4120 2993 4154 3027
rect 4188 2993 4222 3027
rect 4256 2993 4290 3027
rect 4324 2993 4358 3027
rect 4392 2993 4426 3027
rect 4460 2993 4494 3027
rect 4528 2993 4562 3027
rect 4596 2993 4630 3027
rect 4664 2993 4698 3027
rect 4732 2993 4766 3027
rect 4800 2993 4834 3027
rect 4868 2993 4902 3027
rect 4936 2993 4970 3027
rect 5004 2993 5038 3027
rect 5072 2993 5106 3027
rect 5140 2993 5174 3027
rect 5208 2993 5242 3027
rect 5276 2993 5310 3027
rect 5344 2993 5378 3027
rect 5412 2993 5446 3027
rect 5480 2993 5514 3027
rect 5548 2993 5582 3027
rect 5616 2993 5650 3027
rect 5684 2993 5718 3027
rect 5752 2993 5786 3027
rect 5820 2993 5907 3027
rect -557 2938 -523 2993
rect -557 2870 -523 2904
rect -557 2802 -523 2836
rect -557 2734 -523 2768
rect -557 2666 -523 2700
rect -557 2598 -523 2632
rect 5873 2938 5907 2993
rect 5873 2870 5907 2904
rect 5873 2802 5907 2836
rect 5873 2734 5907 2768
rect 5873 2666 5907 2700
rect -557 2530 -523 2564
rect -557 2462 -523 2496
rect -557 2394 -523 2428
rect 5570 2572 5680 2610
rect 5570 2538 5608 2572
rect 5642 2538 5680 2572
rect 5570 2482 5680 2538
rect 5570 2448 5608 2482
rect 5642 2448 5680 2482
rect 5570 2420 5680 2448
rect 5873 2598 5907 2632
rect 5873 2530 5907 2564
rect 5873 2462 5907 2496
rect -557 2326 -523 2360
rect -557 2258 -523 2292
rect -557 2190 -523 2224
rect -557 2122 -523 2156
rect -557 2054 -523 2088
rect -557 1986 -523 2020
rect -557 1918 -523 1952
rect -557 1850 -523 1884
rect -557 1782 -523 1816
rect -557 1714 -523 1748
rect -557 1646 -523 1680
rect -557 1578 -523 1612
rect -557 1510 -523 1544
rect -557 1442 -523 1476
rect -557 1374 -523 1408
rect -557 1306 -523 1340
rect -557 1238 -523 1272
rect -557 1170 -523 1204
rect -557 1102 -523 1136
rect -557 1034 -523 1068
rect -557 966 -523 1000
rect -557 898 -523 932
rect -557 830 -523 864
rect -557 762 -523 796
rect -557 694 -523 728
rect -557 626 -523 660
rect -557 558 -523 592
rect -557 490 -523 524
rect -557 422 -523 456
rect -557 354 -523 388
rect -557 286 -523 320
rect -557 218 -523 252
rect -557 150 -523 184
rect -557 82 -523 116
rect -557 14 -523 48
rect -557 -54 -523 -20
rect -557 -122 -523 -88
rect -557 -190 -523 -156
rect -557 -258 -523 -224
rect -557 -326 -523 -292
rect -557 -394 -523 -360
rect -557 -462 -523 -428
rect -557 -530 -523 -496
rect -557 -598 -523 -564
rect -557 -666 -523 -632
rect -557 -734 -523 -700
rect -557 -802 -523 -768
rect -557 -870 -523 -836
rect -557 -938 -523 -904
rect -557 -1006 -523 -972
rect -557 -1074 -523 -1040
rect -557 -1142 -523 -1108
rect -557 -1210 -523 -1176
rect -557 -1278 -523 -1244
rect -557 -1346 -523 -1312
rect -557 -1414 -523 -1380
rect -557 -1482 -523 -1448
rect -557 -1550 -523 -1516
rect -557 -1618 -523 -1584
rect -557 -1686 -523 -1652
rect -557 -1754 -523 -1720
rect -557 -1822 -523 -1788
rect -557 -1890 -523 -1856
rect -557 -1958 -523 -1924
rect -557 -2026 -523 -1992
rect -557 -2094 -523 -2060
rect -557 -2162 -523 -2128
rect -557 -2230 -523 -2196
rect -557 -2298 -523 -2264
rect -557 -2366 -523 -2332
rect -557 -2434 -523 -2400
rect 5873 2394 5907 2428
rect 5873 2326 5907 2360
rect 5873 2258 5907 2292
rect 5873 2190 5907 2224
rect 5873 2122 5907 2156
rect 5873 2054 5907 2088
rect 5873 1986 5907 2020
rect 5873 1918 5907 1952
rect 5873 1850 5907 1884
rect 5873 1782 5907 1816
rect 5873 1714 5907 1748
rect 5873 1646 5907 1680
rect 5873 1578 5907 1612
rect 5873 1510 5907 1544
rect 5873 1442 5907 1476
rect 5873 1374 5907 1408
rect 5873 1306 5907 1340
rect 5873 1238 5907 1272
rect 5873 1170 5907 1204
rect 5873 1102 5907 1136
rect 5873 1034 5907 1068
rect 5873 966 5907 1000
rect 5873 898 5907 932
rect 5873 830 5907 864
rect 5873 762 5907 796
rect 5873 694 5907 728
rect 5873 626 5907 660
rect 5873 558 5907 592
rect 5873 490 5907 524
rect 5873 422 5907 456
rect 5873 354 5907 388
rect 5873 286 5907 320
rect 5873 218 5907 252
rect 5873 150 5907 184
rect 5873 82 5907 116
rect 5873 14 5907 48
rect 5873 -54 5907 -20
rect 5873 -122 5907 -88
rect 5873 -190 5907 -156
rect 5873 -258 5907 -224
rect 5873 -326 5907 -292
rect 5873 -394 5907 -360
rect 5873 -462 5907 -428
rect 5873 -530 5907 -496
rect 5873 -598 5907 -564
rect 5873 -666 5907 -632
rect 5873 -734 5907 -700
rect 5873 -802 5907 -768
rect 5873 -870 5907 -836
rect 5873 -938 5907 -904
rect 5873 -1006 5907 -972
rect 5873 -1074 5907 -1040
rect 5873 -1142 5907 -1108
rect 5873 -1210 5907 -1176
rect 5873 -1278 5907 -1244
rect 5873 -1346 5907 -1312
rect 5873 -1414 5907 -1380
rect 5873 -1482 5907 -1448
rect 5873 -1550 5907 -1516
rect 5873 -1618 5907 -1584
rect 5873 -1686 5907 -1652
rect 5873 -1754 5907 -1720
rect 5873 -1822 5907 -1788
rect 5873 -1890 5907 -1856
rect 5873 -1958 5907 -1924
rect 5873 -2026 5907 -1992
rect 5873 -2094 5907 -2060
rect 5873 -2162 5907 -2128
rect 5873 -2230 5907 -2196
rect 5873 -2298 5907 -2264
rect 5873 -2366 5907 -2332
rect 5873 -2434 5907 -2400
rect -557 -2502 -523 -2468
rect -557 -2570 -523 -2536
rect -557 -2638 -523 -2604
rect -370 -2498 -260 -2460
rect -370 -2532 -332 -2498
rect -298 -2532 -260 -2498
rect -370 -2588 -260 -2532
rect -370 -2622 -332 -2588
rect -298 -2622 -260 -2588
rect -370 -2650 -260 -2622
rect 5873 -2502 5907 -2468
rect 5873 -2570 5907 -2536
rect 5873 -2638 5907 -2604
rect -557 -2706 -523 -2672
rect -557 -2774 -523 -2740
rect -557 -2863 -523 -2808
rect 5873 -2706 5907 -2672
rect 5873 -2774 5907 -2740
rect 5873 -2863 5907 -2808
rect -557 -2897 -470 -2863
rect -436 -2897 -402 -2863
rect -368 -2897 -334 -2863
rect -300 -2897 -266 -2863
rect -232 -2897 -198 -2863
rect -164 -2897 -130 -2863
rect -96 -2897 -62 -2863
rect -28 -2897 6 -2863
rect 40 -2897 74 -2863
rect 108 -2897 142 -2863
rect 176 -2897 210 -2863
rect 244 -2897 278 -2863
rect 312 -2897 346 -2863
rect 380 -2897 414 -2863
rect 448 -2897 482 -2863
rect 516 -2897 550 -2863
rect 584 -2897 618 -2863
rect 652 -2897 686 -2863
rect 720 -2897 754 -2863
rect 788 -2897 822 -2863
rect 856 -2897 890 -2863
rect 924 -2897 958 -2863
rect 992 -2897 1026 -2863
rect 1060 -2897 1094 -2863
rect 1128 -2897 1162 -2863
rect 1196 -2897 1230 -2863
rect 1264 -2897 1298 -2863
rect 1332 -2897 1366 -2863
rect 1400 -2897 1434 -2863
rect 1468 -2897 1502 -2863
rect 1536 -2897 1570 -2863
rect 1604 -2897 1638 -2863
rect 1672 -2897 1706 -2863
rect 1740 -2897 1774 -2863
rect 1808 -2897 1842 -2863
rect 1876 -2897 1910 -2863
rect 1944 -2897 1978 -2863
rect 2012 -2897 2046 -2863
rect 2080 -2897 2114 -2863
rect 2148 -2897 2182 -2863
rect 2216 -2897 2250 -2863
rect 2284 -2897 2318 -2863
rect 2352 -2897 2386 -2863
rect 2420 -2897 2454 -2863
rect 2488 -2897 2522 -2863
rect 2556 -2897 2590 -2863
rect 2624 -2897 2658 -2863
rect 2692 -2897 2726 -2863
rect 2760 -2897 2794 -2863
rect 2828 -2897 2862 -2863
rect 2896 -2897 2930 -2863
rect 2964 -2897 2998 -2863
rect 3032 -2897 3066 -2863
rect 3100 -2897 3134 -2863
rect 3168 -2897 3202 -2863
rect 3236 -2897 3270 -2863
rect 3304 -2897 3338 -2863
rect 3372 -2897 3406 -2863
rect 3440 -2897 3474 -2863
rect 3508 -2897 3542 -2863
rect 3576 -2897 3610 -2863
rect 3644 -2897 3678 -2863
rect 3712 -2897 3746 -2863
rect 3780 -2897 3814 -2863
rect 3848 -2897 3882 -2863
rect 3916 -2897 3950 -2863
rect 3984 -2897 4018 -2863
rect 4052 -2897 4086 -2863
rect 4120 -2897 4154 -2863
rect 4188 -2897 4222 -2863
rect 4256 -2897 4290 -2863
rect 4324 -2897 4358 -2863
rect 4392 -2897 4426 -2863
rect 4460 -2897 4494 -2863
rect 4528 -2897 4562 -2863
rect 4596 -2897 4630 -2863
rect 4664 -2897 4698 -2863
rect 4732 -2897 4766 -2863
rect 4800 -2897 4834 -2863
rect 4868 -2897 4902 -2863
rect 4936 -2897 4970 -2863
rect 5004 -2897 5038 -2863
rect 5072 -2897 5106 -2863
rect 5140 -2897 5174 -2863
rect 5208 -2897 5242 -2863
rect 5276 -2897 5310 -2863
rect 5344 -2897 5378 -2863
rect 5412 -2897 5446 -2863
rect 5480 -2897 5514 -2863
rect 5548 -2897 5582 -2863
rect 5616 -2897 5650 -2863
rect 5684 -2897 5718 -2863
rect 5752 -2897 5786 -2863
rect 5820 -2897 5907 -2863
<< psubdiffcont >>
rect -470 2993 -436 3027
rect -402 2993 -368 3027
rect -334 2993 -300 3027
rect -266 2993 -232 3027
rect -198 2993 -164 3027
rect -130 2993 -96 3027
rect -62 2993 -28 3027
rect 6 2993 40 3027
rect 74 2993 108 3027
rect 142 2993 176 3027
rect 210 2993 244 3027
rect 278 2993 312 3027
rect 346 2993 380 3027
rect 414 2993 448 3027
rect 482 2993 516 3027
rect 550 2993 584 3027
rect 618 2993 652 3027
rect 686 2993 720 3027
rect 754 2993 788 3027
rect 822 2993 856 3027
rect 890 2993 924 3027
rect 958 2993 992 3027
rect 1026 2993 1060 3027
rect 1094 2993 1128 3027
rect 1162 2993 1196 3027
rect 1230 2993 1264 3027
rect 1298 2993 1332 3027
rect 1366 2993 1400 3027
rect 1434 2993 1468 3027
rect 1502 2993 1536 3027
rect 1570 2993 1604 3027
rect 1638 2993 1672 3027
rect 1706 2993 1740 3027
rect 1774 2993 1808 3027
rect 1842 2993 1876 3027
rect 1910 2993 1944 3027
rect 1978 2993 2012 3027
rect 2046 2993 2080 3027
rect 2114 2993 2148 3027
rect 2182 2993 2216 3027
rect 2250 2993 2284 3027
rect 2318 2993 2352 3027
rect 2386 2993 2420 3027
rect 2454 2993 2488 3027
rect 2522 2993 2556 3027
rect 2590 2993 2624 3027
rect 2658 2993 2692 3027
rect 2726 2993 2760 3027
rect 2794 2993 2828 3027
rect 2862 2993 2896 3027
rect 2930 2993 2964 3027
rect 2998 2993 3032 3027
rect 3066 2993 3100 3027
rect 3134 2993 3168 3027
rect 3202 2993 3236 3027
rect 3270 2993 3304 3027
rect 3338 2993 3372 3027
rect 3406 2993 3440 3027
rect 3474 2993 3508 3027
rect 3542 2993 3576 3027
rect 3610 2993 3644 3027
rect 3678 2993 3712 3027
rect 3746 2993 3780 3027
rect 3814 2993 3848 3027
rect 3882 2993 3916 3027
rect 3950 2993 3984 3027
rect 4018 2993 4052 3027
rect 4086 2993 4120 3027
rect 4154 2993 4188 3027
rect 4222 2993 4256 3027
rect 4290 2993 4324 3027
rect 4358 2993 4392 3027
rect 4426 2993 4460 3027
rect 4494 2993 4528 3027
rect 4562 2993 4596 3027
rect 4630 2993 4664 3027
rect 4698 2993 4732 3027
rect 4766 2993 4800 3027
rect 4834 2993 4868 3027
rect 4902 2993 4936 3027
rect 4970 2993 5004 3027
rect 5038 2993 5072 3027
rect 5106 2993 5140 3027
rect 5174 2993 5208 3027
rect 5242 2993 5276 3027
rect 5310 2993 5344 3027
rect 5378 2993 5412 3027
rect 5446 2993 5480 3027
rect 5514 2993 5548 3027
rect 5582 2993 5616 3027
rect 5650 2993 5684 3027
rect 5718 2993 5752 3027
rect 5786 2993 5820 3027
rect -557 2904 -523 2938
rect -557 2836 -523 2870
rect -557 2768 -523 2802
rect -557 2700 -523 2734
rect -557 2632 -523 2666
rect 5873 2904 5907 2938
rect 5873 2836 5907 2870
rect 5873 2768 5907 2802
rect 5873 2700 5907 2734
rect 5873 2632 5907 2666
rect -557 2564 -523 2598
rect -557 2496 -523 2530
rect -557 2428 -523 2462
rect 5608 2538 5642 2572
rect 5608 2448 5642 2482
rect 5873 2564 5907 2598
rect 5873 2496 5907 2530
rect 5873 2428 5907 2462
rect -557 2360 -523 2394
rect -557 2292 -523 2326
rect -557 2224 -523 2258
rect -557 2156 -523 2190
rect -557 2088 -523 2122
rect -557 2020 -523 2054
rect -557 1952 -523 1986
rect -557 1884 -523 1918
rect -557 1816 -523 1850
rect -557 1748 -523 1782
rect -557 1680 -523 1714
rect -557 1612 -523 1646
rect -557 1544 -523 1578
rect -557 1476 -523 1510
rect -557 1408 -523 1442
rect -557 1340 -523 1374
rect -557 1272 -523 1306
rect -557 1204 -523 1238
rect -557 1136 -523 1170
rect -557 1068 -523 1102
rect -557 1000 -523 1034
rect -557 932 -523 966
rect -557 864 -523 898
rect -557 796 -523 830
rect -557 728 -523 762
rect -557 660 -523 694
rect -557 592 -523 626
rect -557 524 -523 558
rect -557 456 -523 490
rect -557 388 -523 422
rect -557 320 -523 354
rect -557 252 -523 286
rect -557 184 -523 218
rect -557 116 -523 150
rect -557 48 -523 82
rect -557 -20 -523 14
rect -557 -88 -523 -54
rect -557 -156 -523 -122
rect -557 -224 -523 -190
rect -557 -292 -523 -258
rect -557 -360 -523 -326
rect -557 -428 -523 -394
rect -557 -496 -523 -462
rect -557 -564 -523 -530
rect -557 -632 -523 -598
rect -557 -700 -523 -666
rect -557 -768 -523 -734
rect -557 -836 -523 -802
rect -557 -904 -523 -870
rect -557 -972 -523 -938
rect -557 -1040 -523 -1006
rect -557 -1108 -523 -1074
rect -557 -1176 -523 -1142
rect -557 -1244 -523 -1210
rect -557 -1312 -523 -1278
rect -557 -1380 -523 -1346
rect -557 -1448 -523 -1414
rect -557 -1516 -523 -1482
rect -557 -1584 -523 -1550
rect -557 -1652 -523 -1618
rect -557 -1720 -523 -1686
rect -557 -1788 -523 -1754
rect -557 -1856 -523 -1822
rect -557 -1924 -523 -1890
rect -557 -1992 -523 -1958
rect -557 -2060 -523 -2026
rect -557 -2128 -523 -2094
rect -557 -2196 -523 -2162
rect -557 -2264 -523 -2230
rect -557 -2332 -523 -2298
rect -557 -2400 -523 -2366
rect -557 -2468 -523 -2434
rect 5873 2360 5907 2394
rect 5873 2292 5907 2326
rect 5873 2224 5907 2258
rect 5873 2156 5907 2190
rect 5873 2088 5907 2122
rect 5873 2020 5907 2054
rect 5873 1952 5907 1986
rect 5873 1884 5907 1918
rect 5873 1816 5907 1850
rect 5873 1748 5907 1782
rect 5873 1680 5907 1714
rect 5873 1612 5907 1646
rect 5873 1544 5907 1578
rect 5873 1476 5907 1510
rect 5873 1408 5907 1442
rect 5873 1340 5907 1374
rect 5873 1272 5907 1306
rect 5873 1204 5907 1238
rect 5873 1136 5907 1170
rect 5873 1068 5907 1102
rect 5873 1000 5907 1034
rect 5873 932 5907 966
rect 5873 864 5907 898
rect 5873 796 5907 830
rect 5873 728 5907 762
rect 5873 660 5907 694
rect 5873 592 5907 626
rect 5873 524 5907 558
rect 5873 456 5907 490
rect 5873 388 5907 422
rect 5873 320 5907 354
rect 5873 252 5907 286
rect 5873 184 5907 218
rect 5873 116 5907 150
rect 5873 48 5907 82
rect 5873 -20 5907 14
rect 5873 -88 5907 -54
rect 5873 -156 5907 -122
rect 5873 -224 5907 -190
rect 5873 -292 5907 -258
rect 5873 -360 5907 -326
rect 5873 -428 5907 -394
rect 5873 -496 5907 -462
rect 5873 -564 5907 -530
rect 5873 -632 5907 -598
rect 5873 -700 5907 -666
rect 5873 -768 5907 -734
rect 5873 -836 5907 -802
rect 5873 -904 5907 -870
rect 5873 -972 5907 -938
rect 5873 -1040 5907 -1006
rect 5873 -1108 5907 -1074
rect 5873 -1176 5907 -1142
rect 5873 -1244 5907 -1210
rect 5873 -1312 5907 -1278
rect 5873 -1380 5907 -1346
rect 5873 -1448 5907 -1414
rect 5873 -1516 5907 -1482
rect 5873 -1584 5907 -1550
rect 5873 -1652 5907 -1618
rect 5873 -1720 5907 -1686
rect 5873 -1788 5907 -1754
rect 5873 -1856 5907 -1822
rect 5873 -1924 5907 -1890
rect 5873 -1992 5907 -1958
rect 5873 -2060 5907 -2026
rect 5873 -2128 5907 -2094
rect 5873 -2196 5907 -2162
rect 5873 -2264 5907 -2230
rect 5873 -2332 5907 -2298
rect 5873 -2400 5907 -2366
rect -557 -2536 -523 -2502
rect -557 -2604 -523 -2570
rect -557 -2672 -523 -2638
rect -332 -2532 -298 -2498
rect -332 -2622 -298 -2588
rect 5873 -2468 5907 -2434
rect 5873 -2536 5907 -2502
rect 5873 -2604 5907 -2570
rect -557 -2740 -523 -2706
rect -557 -2808 -523 -2774
rect 5873 -2672 5907 -2638
rect 5873 -2740 5907 -2706
rect 5873 -2808 5907 -2774
rect -470 -2897 -436 -2863
rect -402 -2897 -368 -2863
rect -334 -2897 -300 -2863
rect -266 -2897 -232 -2863
rect -198 -2897 -164 -2863
rect -130 -2897 -96 -2863
rect -62 -2897 -28 -2863
rect 6 -2897 40 -2863
rect 74 -2897 108 -2863
rect 142 -2897 176 -2863
rect 210 -2897 244 -2863
rect 278 -2897 312 -2863
rect 346 -2897 380 -2863
rect 414 -2897 448 -2863
rect 482 -2897 516 -2863
rect 550 -2897 584 -2863
rect 618 -2897 652 -2863
rect 686 -2897 720 -2863
rect 754 -2897 788 -2863
rect 822 -2897 856 -2863
rect 890 -2897 924 -2863
rect 958 -2897 992 -2863
rect 1026 -2897 1060 -2863
rect 1094 -2897 1128 -2863
rect 1162 -2897 1196 -2863
rect 1230 -2897 1264 -2863
rect 1298 -2897 1332 -2863
rect 1366 -2897 1400 -2863
rect 1434 -2897 1468 -2863
rect 1502 -2897 1536 -2863
rect 1570 -2897 1604 -2863
rect 1638 -2897 1672 -2863
rect 1706 -2897 1740 -2863
rect 1774 -2897 1808 -2863
rect 1842 -2897 1876 -2863
rect 1910 -2897 1944 -2863
rect 1978 -2897 2012 -2863
rect 2046 -2897 2080 -2863
rect 2114 -2897 2148 -2863
rect 2182 -2897 2216 -2863
rect 2250 -2897 2284 -2863
rect 2318 -2897 2352 -2863
rect 2386 -2897 2420 -2863
rect 2454 -2897 2488 -2863
rect 2522 -2897 2556 -2863
rect 2590 -2897 2624 -2863
rect 2658 -2897 2692 -2863
rect 2726 -2897 2760 -2863
rect 2794 -2897 2828 -2863
rect 2862 -2897 2896 -2863
rect 2930 -2897 2964 -2863
rect 2998 -2897 3032 -2863
rect 3066 -2897 3100 -2863
rect 3134 -2897 3168 -2863
rect 3202 -2897 3236 -2863
rect 3270 -2897 3304 -2863
rect 3338 -2897 3372 -2863
rect 3406 -2897 3440 -2863
rect 3474 -2897 3508 -2863
rect 3542 -2897 3576 -2863
rect 3610 -2897 3644 -2863
rect 3678 -2897 3712 -2863
rect 3746 -2897 3780 -2863
rect 3814 -2897 3848 -2863
rect 3882 -2897 3916 -2863
rect 3950 -2897 3984 -2863
rect 4018 -2897 4052 -2863
rect 4086 -2897 4120 -2863
rect 4154 -2897 4188 -2863
rect 4222 -2897 4256 -2863
rect 4290 -2897 4324 -2863
rect 4358 -2897 4392 -2863
rect 4426 -2897 4460 -2863
rect 4494 -2897 4528 -2863
rect 4562 -2897 4596 -2863
rect 4630 -2897 4664 -2863
rect 4698 -2897 4732 -2863
rect 4766 -2897 4800 -2863
rect 4834 -2897 4868 -2863
rect 4902 -2897 4936 -2863
rect 4970 -2897 5004 -2863
rect 5038 -2897 5072 -2863
rect 5106 -2897 5140 -2863
rect 5174 -2897 5208 -2863
rect 5242 -2897 5276 -2863
rect 5310 -2897 5344 -2863
rect 5378 -2897 5412 -2863
rect 5446 -2897 5480 -2863
rect 5514 -2897 5548 -2863
rect 5582 -2897 5616 -2863
rect 5650 -2897 5684 -2863
rect 5718 -2897 5752 -2863
rect 5786 -2897 5820 -2863
<< locali >>
rect -557 2993 -470 3027
rect -436 2993 -402 3027
rect -368 2993 -334 3027
rect -300 2993 -266 3027
rect -232 2993 -198 3027
rect -164 2993 -130 3027
rect -96 2993 -62 3027
rect -28 2993 6 3027
rect 40 2993 74 3027
rect 108 2993 142 3027
rect 176 2993 210 3027
rect 244 2993 278 3027
rect 312 2993 346 3027
rect 380 2993 414 3027
rect 448 2993 482 3027
rect 516 2993 550 3027
rect 584 2993 618 3027
rect 652 2993 686 3027
rect 720 2993 754 3027
rect 788 2993 822 3027
rect 856 2993 890 3027
rect 924 2993 958 3027
rect 992 2993 1026 3027
rect 1060 2993 1094 3027
rect 1128 2993 1162 3027
rect 1196 2993 1230 3027
rect 1264 2993 1298 3027
rect 1332 2993 1366 3027
rect 1400 2993 1434 3027
rect 1468 2993 1502 3027
rect 1536 2993 1570 3027
rect 1604 2993 1638 3027
rect 1672 2993 1706 3027
rect 1740 2993 1774 3027
rect 1808 2993 1842 3027
rect 1876 2993 1910 3027
rect 1944 2993 1978 3027
rect 2012 2993 2046 3027
rect 2080 2993 2114 3027
rect 2148 2993 2182 3027
rect 2216 2993 2250 3027
rect 2284 2993 2318 3027
rect 2352 2993 2386 3027
rect 2420 2993 2454 3027
rect 2488 2993 2522 3027
rect 2556 2993 2590 3027
rect 2624 2993 2658 3027
rect 2692 2993 2726 3027
rect 2760 2993 2794 3027
rect 2828 2993 2862 3027
rect 2896 2993 2930 3027
rect 2964 2993 2998 3027
rect 3032 2993 3066 3027
rect 3100 2993 3134 3027
rect 3168 2993 3202 3027
rect 3236 2993 3270 3027
rect 3304 2993 3338 3027
rect 3372 2993 3406 3027
rect 3440 2993 3474 3027
rect 3508 2993 3542 3027
rect 3576 2993 3610 3027
rect 3644 2993 3678 3027
rect 3712 2993 3746 3027
rect 3780 2993 3814 3027
rect 3848 2993 3882 3027
rect 3916 2993 3950 3027
rect 3984 2993 4018 3027
rect 4052 2993 4086 3027
rect 4120 2993 4154 3027
rect 4188 2993 4222 3027
rect 4256 2993 4290 3027
rect 4324 2993 4358 3027
rect 4392 2993 4426 3027
rect 4460 2993 4494 3027
rect 4528 2993 4562 3027
rect 4596 2993 4630 3027
rect 4664 2993 4698 3027
rect 4732 2993 4766 3027
rect 4800 2993 4834 3027
rect 4868 2993 4902 3027
rect 4936 2993 4970 3027
rect 5004 2993 5038 3027
rect 5072 2993 5106 3027
rect 5140 2993 5174 3027
rect 5208 2993 5242 3027
rect 5276 2993 5310 3027
rect 5344 2993 5378 3027
rect 5412 2993 5446 3027
rect 5480 2993 5514 3027
rect 5548 2993 5582 3027
rect 5616 2993 5650 3027
rect 5684 2993 5718 3027
rect 5752 2993 5786 3027
rect 5820 2993 5907 3027
rect -557 2938 -523 2993
rect -557 2870 -523 2904
rect -557 2802 -523 2836
rect -557 2734 -523 2768
rect -557 2666 -523 2700
rect -557 2598 -523 2632
rect 5873 2938 5907 2993
rect 5873 2870 5907 2904
rect 5873 2802 5907 2836
rect 5873 2734 5907 2768
rect 5873 2666 5907 2700
rect -557 2530 -523 2564
rect -557 2462 -523 2496
rect -557 2394 -523 2428
rect 5570 2572 5680 2610
rect 5570 2538 5608 2572
rect 5642 2538 5680 2572
rect 5570 2482 5680 2538
rect 5570 2448 5608 2482
rect 5642 2448 5680 2482
rect 5570 2420 5680 2448
rect 5873 2598 5907 2632
rect 5873 2530 5907 2564
rect 5873 2462 5907 2496
rect -557 2326 -523 2360
rect -557 2258 -523 2292
rect -557 2190 -523 2224
rect -557 2122 -523 2156
rect -557 2054 -523 2088
rect -557 1986 -523 2020
rect -557 1918 -523 1952
rect -557 1850 -523 1884
rect -557 1782 -523 1816
rect -557 1714 -523 1748
rect -557 1646 -523 1680
rect -557 1578 -523 1612
rect -557 1510 -523 1544
rect -557 1442 -523 1476
rect -557 1374 -523 1408
rect -557 1306 -523 1340
rect -557 1238 -523 1272
rect -557 1170 -523 1204
rect -557 1102 -523 1136
rect -557 1034 -523 1068
rect -557 966 -523 1000
rect -557 898 -523 932
rect -557 830 -523 864
rect -557 762 -523 796
rect -557 694 -523 728
rect -557 626 -523 660
rect -557 558 -523 592
rect -557 490 -523 524
rect -557 422 -523 456
rect -557 354 -523 388
rect -557 286 -523 320
rect -557 218 -523 252
rect -557 150 -523 184
rect -557 82 -523 116
rect -557 14 -523 48
rect -557 -54 -523 -20
rect -557 -122 -523 -88
rect -557 -190 -523 -156
rect -557 -258 -523 -224
rect -557 -326 -523 -292
rect -557 -394 -523 -360
rect -557 -462 -523 -428
rect -557 -530 -523 -496
rect -557 -598 -523 -564
rect -557 -666 -523 -632
rect -557 -734 -523 -700
rect -557 -802 -523 -768
rect -557 -870 -523 -836
rect -557 -938 -523 -904
rect -557 -1006 -523 -972
rect -557 -1074 -523 -1040
rect -557 -1142 -523 -1108
rect -557 -1210 -523 -1176
rect -557 -1278 -523 -1244
rect -557 -1346 -523 -1312
rect -557 -1414 -523 -1380
rect -557 -1482 -523 -1448
rect -557 -1550 -523 -1516
rect -557 -1618 -523 -1584
rect -557 -1686 -523 -1652
rect -557 -1754 -523 -1720
rect -557 -1822 -523 -1788
rect -557 -1890 -523 -1856
rect -557 -1958 -523 -1924
rect -557 -2026 -523 -1992
rect -557 -2094 -523 -2060
rect -557 -2162 -523 -2128
rect -557 -2230 -523 -2196
rect -557 -2298 -523 -2264
rect -557 -2366 -523 -2332
rect -557 -2434 -523 -2400
rect 5873 2394 5907 2428
rect 5873 2326 5907 2360
rect 5873 2258 5907 2292
rect 5873 2190 5907 2224
rect 5873 2122 5907 2156
rect 5873 2054 5907 2088
rect 5873 1986 5907 2020
rect 5873 1918 5907 1952
rect 5873 1850 5907 1884
rect 5873 1782 5907 1816
rect 5873 1714 5907 1748
rect 5873 1646 5907 1680
rect 5873 1578 5907 1612
rect 5873 1510 5907 1544
rect 5873 1442 5907 1476
rect 5873 1374 5907 1408
rect 5873 1306 5907 1340
rect 5873 1238 5907 1272
rect 5873 1170 5907 1204
rect 5873 1102 5907 1136
rect 5873 1034 5907 1068
rect 5873 966 5907 1000
rect 5873 898 5907 932
rect 5873 830 5907 864
rect 5873 762 5907 796
rect 5873 694 5907 728
rect 5873 626 5907 660
rect 5873 558 5907 592
rect 5873 490 5907 524
rect 5873 422 5907 456
rect 5873 354 5907 388
rect 5873 286 5907 320
rect 5873 218 5907 252
rect 5873 150 5907 184
rect 5873 82 5907 116
rect 5873 14 5907 48
rect 5873 -54 5907 -20
rect 5873 -122 5907 -88
rect 5873 -190 5907 -156
rect 5873 -258 5907 -224
rect 5873 -326 5907 -292
rect 5873 -394 5907 -360
rect 5873 -462 5907 -428
rect 5873 -530 5907 -496
rect 5873 -598 5907 -564
rect 5873 -666 5907 -632
rect 5873 -734 5907 -700
rect 5873 -802 5907 -768
rect 5873 -870 5907 -836
rect 5873 -938 5907 -904
rect 5873 -1006 5907 -972
rect 5873 -1074 5907 -1040
rect 5873 -1142 5907 -1108
rect 5873 -1210 5907 -1176
rect 5873 -1278 5907 -1244
rect 5873 -1346 5907 -1312
rect 5873 -1414 5907 -1380
rect 5873 -1482 5907 -1448
rect 5873 -1550 5907 -1516
rect 5873 -1618 5907 -1584
rect 5873 -1686 5907 -1652
rect 5873 -1754 5907 -1720
rect 5873 -1822 5907 -1788
rect 5873 -1890 5907 -1856
rect 5873 -1958 5907 -1924
rect 5873 -2026 5907 -1992
rect 5873 -2094 5907 -2060
rect 5873 -2162 5907 -2128
rect 5873 -2230 5907 -2196
rect 5873 -2298 5907 -2264
rect 5873 -2366 5907 -2332
rect 5873 -2434 5907 -2400
rect -557 -2502 -523 -2468
rect -557 -2570 -523 -2536
rect -557 -2638 -523 -2604
rect -370 -2498 -260 -2460
rect -370 -2532 -332 -2498
rect -298 -2532 -260 -2498
rect -370 -2588 -260 -2532
rect -370 -2622 -332 -2588
rect -298 -2622 -260 -2588
rect -370 -2650 -260 -2622
rect 5873 -2502 5907 -2468
rect 5873 -2570 5907 -2536
rect 5873 -2638 5907 -2604
rect -557 -2706 -523 -2672
rect -557 -2774 -523 -2740
rect -557 -2863 -523 -2808
rect 5873 -2706 5907 -2672
rect 5873 -2774 5907 -2740
rect 5873 -2863 5907 -2808
rect -557 -2897 -470 -2863
rect -436 -2897 -402 -2863
rect -368 -2897 -334 -2863
rect -300 -2897 -266 -2863
rect -232 -2897 -198 -2863
rect -164 -2897 -130 -2863
rect -96 -2897 -62 -2863
rect -28 -2897 6 -2863
rect 40 -2897 74 -2863
rect 108 -2897 142 -2863
rect 176 -2897 210 -2863
rect 244 -2897 278 -2863
rect 312 -2897 346 -2863
rect 380 -2897 414 -2863
rect 448 -2897 482 -2863
rect 516 -2897 550 -2863
rect 584 -2897 618 -2863
rect 652 -2897 686 -2863
rect 720 -2897 754 -2863
rect 788 -2897 822 -2863
rect 856 -2897 890 -2863
rect 924 -2897 958 -2863
rect 992 -2897 1026 -2863
rect 1060 -2897 1094 -2863
rect 1128 -2897 1162 -2863
rect 1196 -2897 1230 -2863
rect 1264 -2897 1298 -2863
rect 1332 -2897 1366 -2863
rect 1400 -2897 1434 -2863
rect 1468 -2897 1502 -2863
rect 1536 -2897 1570 -2863
rect 1604 -2897 1638 -2863
rect 1672 -2897 1706 -2863
rect 1740 -2897 1774 -2863
rect 1808 -2897 1842 -2863
rect 1876 -2897 1910 -2863
rect 1944 -2897 1978 -2863
rect 2012 -2897 2046 -2863
rect 2080 -2897 2114 -2863
rect 2148 -2897 2182 -2863
rect 2216 -2897 2250 -2863
rect 2284 -2897 2318 -2863
rect 2352 -2897 2386 -2863
rect 2420 -2897 2454 -2863
rect 2488 -2897 2522 -2863
rect 2556 -2897 2590 -2863
rect 2624 -2897 2658 -2863
rect 2692 -2897 2726 -2863
rect 2760 -2897 2794 -2863
rect 2828 -2897 2862 -2863
rect 2896 -2897 2930 -2863
rect 2964 -2897 2998 -2863
rect 3032 -2897 3066 -2863
rect 3100 -2897 3134 -2863
rect 3168 -2897 3202 -2863
rect 3236 -2897 3270 -2863
rect 3304 -2897 3338 -2863
rect 3372 -2897 3406 -2863
rect 3440 -2897 3474 -2863
rect 3508 -2897 3542 -2863
rect 3576 -2897 3610 -2863
rect 3644 -2897 3678 -2863
rect 3712 -2897 3746 -2863
rect 3780 -2897 3814 -2863
rect 3848 -2897 3882 -2863
rect 3916 -2897 3950 -2863
rect 3984 -2897 4018 -2863
rect 4052 -2897 4086 -2863
rect 4120 -2897 4154 -2863
rect 4188 -2897 4222 -2863
rect 4256 -2897 4290 -2863
rect 4324 -2897 4358 -2863
rect 4392 -2897 4426 -2863
rect 4460 -2897 4494 -2863
rect 4528 -2897 4562 -2863
rect 4596 -2897 4630 -2863
rect 4664 -2897 4698 -2863
rect 4732 -2897 4766 -2863
rect 4800 -2897 4834 -2863
rect 4868 -2897 4902 -2863
rect 4936 -2897 4970 -2863
rect 5004 -2897 5038 -2863
rect 5072 -2897 5106 -2863
rect 5140 -2897 5174 -2863
rect 5208 -2897 5242 -2863
rect 5276 -2897 5310 -2863
rect 5344 -2897 5378 -2863
rect 5412 -2897 5446 -2863
rect 5480 -2897 5514 -2863
rect 5548 -2897 5582 -2863
rect 5616 -2897 5650 -2863
rect 5684 -2897 5718 -2863
rect 5752 -2897 5786 -2863
rect 5820 -2897 5907 -2863
<< viali >>
rect 5608 2538 5642 2572
rect 5608 2448 5642 2482
rect -332 -2532 -298 -2498
rect -332 -2622 -298 -2588
<< metal1 >>
rect -390 2706 -310 2710
rect -390 2654 -376 2706
rect -324 2654 -310 2706
rect -390 2650 -310 2654
rect -390 2286 -330 2650
rect -200 2572 5690 2630
rect -200 2538 5608 2572
rect 5642 2538 5690 2572
rect -200 2482 5690 2538
rect -200 2448 5608 2482
rect 5642 2448 5690 2482
rect -200 2410 5690 2448
rect -190 2330 -10 2410
rect -390 2234 -386 2286
rect -334 2234 -330 2286
rect -390 2206 -330 2234
rect -390 2154 -386 2206
rect -334 2154 -330 2206
rect -390 2140 -330 2154
rect -300 2296 -140 2300
rect -300 2244 -286 2296
rect -234 2244 -206 2296
rect -154 2244 -140 2296
rect -300 2240 -140 2244
rect -480 46 -420 60
rect -480 -6 -476 46
rect -424 -6 -420 46
rect -480 -34 -420 -6
rect -480 -86 -476 -34
rect -424 -86 -420 -34
rect -480 -2770 -420 -86
rect -390 -44 -330 -30
rect -390 -96 -386 -44
rect -334 -96 -330 -44
rect -390 -124 -330 -96
rect -390 -176 -386 -124
rect -334 -176 -330 -124
rect -390 -2184 -330 -176
rect -390 -2236 -386 -2184
rect -334 -2236 -330 -2184
rect -390 -2264 -330 -2236
rect -390 -2316 -386 -2264
rect -334 -2316 -330 -2264
rect -390 -2330 -330 -2316
rect -300 -2360 -240 2240
rect -110 2210 -10 2330
rect 5270 2210 5440 2410
rect 5470 2296 5630 2300
rect 5470 2244 5484 2296
rect 5536 2244 5564 2296
rect 5616 2244 5630 2296
rect 5470 2240 5630 2244
rect -190 2150 -10 2210
rect 70 2150 250 2210
rect 330 2150 510 2210
rect 590 2206 940 2210
rect 590 2154 604 2206
rect 656 2154 704 2206
rect 756 2154 804 2206
rect 856 2154 940 2206
rect 590 2150 940 2154
rect 1110 2150 1290 2210
rect 1370 2206 1720 2210
rect 1370 2154 1394 2206
rect 1446 2154 1514 2206
rect 1566 2154 1634 2206
rect 1686 2154 1720 2206
rect 1370 2150 1720 2154
rect 1890 2206 1980 2210
rect 1890 2154 1909 2206
rect 1961 2154 1980 2206
rect 1890 2150 1980 2154
rect 2150 2150 2330 2210
rect 2410 2150 2590 2210
rect 2670 2150 2850 2210
rect 2930 2150 3110 2210
rect 3190 2206 3280 2210
rect 3190 2154 3209 2206
rect 3261 2154 3280 2206
rect 3190 2150 3280 2154
rect 3450 2206 3800 2210
rect 3450 2154 3474 2206
rect 3526 2154 3604 2206
rect 3656 2154 3734 2206
rect 3786 2154 3800 2206
rect 3450 2150 3800 2154
rect 3970 2150 4150 2210
rect 4230 2206 4580 2210
rect 4230 2154 4254 2206
rect 4306 2154 4384 2206
rect 4436 2154 4504 2206
rect 4556 2154 4580 2206
rect 4230 2150 4580 2154
rect 4750 2150 4930 2210
rect 5010 2150 5190 2210
rect 5270 2150 5450 2210
rect -70 150 -10 2150
rect 190 2030 250 2150
rect 450 2030 510 2150
rect 1230 2030 1290 2150
rect 2270 2030 2330 2150
rect 2530 2030 2590 2150
rect 2790 2030 2850 2150
rect 3050 2030 3110 2150
rect 4090 2030 4150 2150
rect 4870 2030 4930 2150
rect 5130 2030 5190 2150
rect 170 2016 250 2030
rect 170 1964 184 2016
rect 236 1964 250 2016
rect 170 1926 250 1964
rect 170 1874 184 1926
rect 236 1874 250 1926
rect 170 1860 250 1874
rect 430 2016 510 2030
rect 430 1964 444 2016
rect 496 1964 510 2016
rect 430 1926 510 1964
rect 430 1874 444 1926
rect 496 1874 510 1926
rect 430 1860 510 1874
rect 690 2016 770 2030
rect 690 1964 704 2016
rect 756 1964 770 2016
rect 690 1926 770 1964
rect 690 1874 704 1926
rect 756 1874 770 1926
rect 690 1860 770 1874
rect 950 2016 1030 2030
rect 950 1964 964 2016
rect 1016 1964 1030 2016
rect 950 1926 1030 1964
rect 950 1874 964 1926
rect 1016 1874 1030 1926
rect 950 1860 1030 1874
rect 1210 2016 1290 2030
rect 1210 1964 1224 2016
rect 1276 1964 1290 2016
rect 1210 1926 1290 1964
rect 1210 1874 1224 1926
rect 1276 1874 1290 1926
rect 1210 1860 1290 1874
rect 1470 2016 1550 2030
rect 1470 1964 1484 2016
rect 1536 1964 1550 2016
rect 1470 1926 1550 1964
rect 1470 1874 1484 1926
rect 1536 1874 1550 1926
rect 1470 1860 1550 1874
rect 1730 2016 1810 2030
rect 1730 1964 1744 2016
rect 1796 1964 1810 2016
rect 1730 1926 1810 1964
rect 1730 1874 1744 1926
rect 1796 1874 1810 1926
rect 1730 1860 1810 1874
rect 1990 2016 2070 2030
rect 1990 1964 2004 2016
rect 2056 1964 2070 2016
rect 1990 1926 2070 1964
rect 1990 1874 2004 1926
rect 2056 1874 2070 1926
rect 1990 1860 2070 1874
rect 2250 2016 2330 2030
rect 2250 1964 2264 2016
rect 2316 1964 2330 2016
rect 2250 1926 2330 1964
rect 2250 1874 2264 1926
rect 2316 1874 2330 1926
rect 2250 1860 2330 1874
rect 2510 2016 2590 2030
rect 2510 1964 2524 2016
rect 2576 1964 2590 2016
rect 2510 1926 2590 1964
rect 2510 1874 2524 1926
rect 2576 1874 2590 1926
rect 2510 1860 2590 1874
rect 2770 2016 2850 2030
rect 2770 1964 2784 2016
rect 2836 1964 2850 2016
rect 2770 1926 2850 1964
rect 2770 1874 2784 1926
rect 2836 1874 2850 1926
rect 2770 1860 2850 1874
rect 3030 2016 3110 2030
rect 3030 1964 3044 2016
rect 3096 1964 3110 2016
rect 3030 1926 3110 1964
rect 3030 1874 3044 1926
rect 3096 1874 3110 1926
rect 3030 1860 3110 1874
rect 3290 2016 3370 2030
rect 3290 1964 3304 2016
rect 3356 1964 3370 2016
rect 3290 1926 3370 1964
rect 3290 1874 3304 1926
rect 3356 1874 3370 1926
rect 3290 1860 3370 1874
rect 3550 2016 3630 2030
rect 3550 1964 3564 2016
rect 3616 1964 3630 2016
rect 3550 1926 3630 1964
rect 3550 1874 3564 1926
rect 3616 1874 3630 1926
rect 3550 1860 3630 1874
rect 3810 2016 3890 2030
rect 3810 1964 3824 2016
rect 3876 1964 3890 2016
rect 3810 1926 3890 1964
rect 3810 1874 3824 1926
rect 3876 1874 3890 1926
rect 3810 1860 3890 1874
rect 4070 2016 4150 2030
rect 4070 1964 4084 2016
rect 4136 1964 4150 2016
rect 4070 1926 4150 1964
rect 4070 1874 4084 1926
rect 4136 1874 4150 1926
rect 4070 1860 4150 1874
rect 4330 2016 4410 2030
rect 4330 1964 4344 2016
rect 4396 1964 4410 2016
rect 4330 1926 4410 1964
rect 4330 1874 4344 1926
rect 4396 1874 4410 1926
rect 4330 1860 4410 1874
rect 4590 2016 4670 2030
rect 4590 1964 4604 2016
rect 4656 1964 4670 2016
rect 4590 1926 4670 1964
rect 4590 1874 4604 1926
rect 4656 1874 4670 1926
rect 4590 1860 4670 1874
rect 4850 2016 4930 2030
rect 4850 1964 4864 2016
rect 4916 1964 4930 2016
rect 4850 1926 4930 1964
rect 4850 1874 4864 1926
rect 4916 1874 4930 1926
rect 4850 1860 4930 1874
rect 5110 2016 5190 2030
rect 5110 1964 5124 2016
rect 5176 1964 5190 2016
rect 5110 1926 5190 1964
rect 5110 1874 5124 1926
rect 5176 1874 5190 1926
rect 5110 1860 5190 1874
rect -190 146 160 150
rect -190 94 -171 146
rect -119 94 -41 146
rect 11 94 89 146
rect 141 94 160 146
rect -190 90 160 94
rect -190 -180 -10 90
rect 190 -120 250 1860
rect 330 146 420 150
rect 330 94 349 146
rect 401 94 420 146
rect 330 90 420 94
rect 450 -120 510 1860
rect 590 146 680 150
rect 590 94 609 146
rect 661 94 680 146
rect 590 90 680 94
rect 70 -180 250 -120
rect 330 -180 510 -120
rect 590 -124 680 -120
rect 590 -176 609 -124
rect 661 -176 680 -124
rect 590 -180 680 -176
rect -70 -2180 -10 -180
rect 190 -1890 250 -180
rect 450 -1890 510 -180
rect 710 -1890 770 1860
rect 850 146 940 150
rect 850 94 869 146
rect 921 94 940 146
rect 850 90 940 94
rect 850 -124 940 -120
rect 850 -176 869 -124
rect 921 -176 940 -124
rect 850 -180 940 -176
rect 970 -1890 1030 1860
rect 1110 146 1200 150
rect 1110 94 1129 146
rect 1181 94 1200 146
rect 1110 90 1200 94
rect 1230 -120 1290 1860
rect 1370 146 1460 150
rect 1370 94 1389 146
rect 1441 94 1460 146
rect 1370 90 1460 94
rect 1110 -180 1290 -120
rect 1370 -124 1460 -120
rect 1370 -176 1389 -124
rect 1441 -176 1460 -124
rect 1370 -180 1460 -176
rect 1230 -1890 1290 -180
rect 1490 -1890 1550 1860
rect 1630 146 1720 150
rect 1630 94 1649 146
rect 1701 94 1720 146
rect 1630 90 1720 94
rect 1630 -124 1720 -120
rect 1630 -176 1649 -124
rect 1701 -176 1720 -124
rect 1630 -180 1720 -176
rect 1750 -1890 1810 1860
rect 1890 146 1980 150
rect 1890 94 1909 146
rect 1961 94 1980 146
rect 1890 90 1980 94
rect 1890 -124 1980 -120
rect 1890 -176 1909 -124
rect 1961 -176 1980 -124
rect 1890 -180 1980 -176
rect 2010 -1890 2070 1860
rect 2150 146 2240 150
rect 2150 94 2169 146
rect 2221 94 2240 146
rect 2150 90 2240 94
rect 2270 -120 2330 1860
rect 2410 146 2500 150
rect 2410 94 2429 146
rect 2481 94 2500 146
rect 2410 90 2500 94
rect 2530 -120 2590 1860
rect 2670 146 2760 150
rect 2670 94 2689 146
rect 2741 94 2760 146
rect 2670 90 2760 94
rect 2790 -120 2850 1860
rect 2930 146 3020 150
rect 2930 94 2949 146
rect 3001 94 3020 146
rect 2930 90 3020 94
rect 3050 -120 3110 1860
rect 3190 146 3280 150
rect 3190 94 3209 146
rect 3261 94 3280 146
rect 3190 90 3280 94
rect 2150 -180 2330 -120
rect 2410 -180 2590 -120
rect 2670 -180 2850 -120
rect 2930 -180 3110 -120
rect 3190 -124 3280 -120
rect 3190 -176 3209 -124
rect 3261 -176 3280 -124
rect 3190 -180 3280 -176
rect 2270 -1890 2330 -180
rect 2530 -1890 2590 -180
rect 2790 -1890 2850 -180
rect 3050 -1890 3110 -180
rect 3310 -1890 3370 1860
rect 3450 146 3540 150
rect 3450 94 3469 146
rect 3521 94 3540 146
rect 3450 90 3540 94
rect 3450 -124 3540 -120
rect 3450 -176 3469 -124
rect 3521 -176 3540 -124
rect 3450 -180 3540 -176
rect 3570 -1890 3630 1860
rect 3710 146 3800 150
rect 3710 94 3729 146
rect 3781 94 3800 146
rect 3710 90 3800 94
rect 3710 -124 3800 -120
rect 3710 -176 3729 -124
rect 3781 -176 3800 -124
rect 3710 -180 3800 -176
rect 3830 -1890 3890 1860
rect 3970 146 4060 150
rect 3970 94 3989 146
rect 4041 94 4060 146
rect 3970 90 4060 94
rect 4090 -120 4150 1860
rect 4230 146 4320 150
rect 4230 94 4249 146
rect 4301 94 4320 146
rect 4230 90 4320 94
rect 3970 -180 4150 -120
rect 4230 -124 4320 -120
rect 4230 -176 4249 -124
rect 4301 -176 4320 -124
rect 4230 -180 4320 -176
rect 4090 -1890 4150 -180
rect 4350 -1890 4410 1860
rect 4490 146 4580 150
rect 4490 94 4509 146
rect 4561 94 4580 146
rect 4490 90 4580 94
rect 4490 -124 4580 -120
rect 4490 -176 4509 -124
rect 4561 -176 4580 -124
rect 4490 -180 4580 -176
rect 4610 -1890 4670 1860
rect 4750 146 4840 150
rect 4750 94 4769 146
rect 4821 94 4840 146
rect 4750 90 4840 94
rect 4870 -120 4930 1860
rect 5010 146 5100 150
rect 5010 94 5029 146
rect 5081 94 5100 146
rect 5010 90 5100 94
rect 5130 -120 5190 1860
rect 5390 150 5450 2150
rect 4750 -180 4930 -120
rect 5010 -180 5190 -120
rect 5240 146 5450 150
rect 5240 94 5254 146
rect 5306 94 5334 146
rect 5386 94 5450 146
rect 5240 90 5450 94
rect 5240 -120 5350 90
rect 5380 -34 5540 -30
rect 5380 -86 5394 -34
rect 5446 -86 5474 -34
rect 5526 -86 5540 -34
rect 5380 -90 5540 -86
rect 5240 -180 5450 -120
rect 4870 -1890 4930 -180
rect 5130 -1890 5190 -180
rect 5390 -2180 5450 -180
rect -190 -2184 5450 -2180
rect -190 -2236 -171 -2184
rect -119 -2236 -81 -2184
rect -29 -2236 89 -2184
rect 141 -2236 349 -2184
rect 401 -2236 609 -2184
rect 661 -2236 869 -2184
rect 921 -2236 1129 -2184
rect 1181 -2236 1389 -2184
rect 1441 -2236 1649 -2184
rect 1701 -2236 1909 -2184
rect 1961 -2236 2169 -2184
rect 2221 -2236 2429 -2184
rect 2481 -2236 2689 -2184
rect 2741 -2236 2949 -2184
rect 3001 -2236 3209 -2184
rect 3261 -2236 3469 -2184
rect 3521 -2236 3729 -2184
rect 3781 -2236 3989 -2184
rect 4041 -2236 4249 -2184
rect 4301 -2236 4509 -2184
rect 4561 -2236 4769 -2184
rect 4821 -2236 5029 -2184
rect 5081 -2236 5144 -2184
rect 5196 -2236 5274 -2184
rect 5326 -2236 5450 -2184
rect -190 -2240 5450 -2236
rect -300 -2364 -140 -2360
rect -300 -2416 -286 -2364
rect -234 -2416 -206 -2364
rect -154 -2416 -140 -2364
rect -300 -2420 -140 -2416
rect -110 -2450 -10 -2240
rect 5480 -2360 5540 -90
rect 5570 -2184 5630 2240
rect 5570 -2236 5574 -2184
rect 5626 -2236 5630 -2184
rect 5570 -2264 5630 -2236
rect 5570 -2316 5574 -2264
rect 5626 -2316 5630 -2264
rect 5570 -2330 5630 -2316
rect 5660 46 5720 60
rect 5660 -6 5664 46
rect 5716 -6 5720 46
rect 5660 -34 5720 -6
rect 5660 -86 5664 -34
rect 5716 -86 5720 -34
rect 5380 -2364 5540 -2360
rect 5380 -2416 5394 -2364
rect 5446 -2416 5474 -2364
rect 5526 -2416 5540 -2364
rect 5380 -2420 5540 -2416
rect -370 -2498 5450 -2450
rect -370 -2532 -332 -2498
rect -298 -2532 5450 -2498
rect -370 -2588 5450 -2532
rect -370 -2622 -332 -2588
rect -298 -2622 5450 -2588
rect -370 -2660 5450 -2622
rect -190 -2670 5450 -2660
rect 5660 -2680 5720 -86
rect 5560 -2684 5720 -2680
rect 5560 -2736 5574 -2684
rect 5626 -2736 5654 -2684
rect 5706 -2736 5720 -2684
rect 5560 -2740 5720 -2736
rect -480 -2774 -320 -2770
rect -480 -2826 -466 -2774
rect -414 -2826 -386 -2774
rect -334 -2826 -320 -2774
rect -480 -2830 -320 -2826
<< via1 >>
rect -376 2654 -324 2706
rect -386 2234 -334 2286
rect -386 2154 -334 2206
rect -286 2244 -234 2296
rect -206 2244 -154 2296
rect -476 -6 -424 46
rect -476 -86 -424 -34
rect -386 -96 -334 -44
rect -386 -176 -334 -124
rect -386 -2236 -334 -2184
rect -386 -2316 -334 -2264
rect 5484 2244 5536 2296
rect 5564 2244 5616 2296
rect 604 2154 656 2206
rect 704 2154 756 2206
rect 804 2154 856 2206
rect 1394 2154 1446 2206
rect 1514 2154 1566 2206
rect 1634 2154 1686 2206
rect 1909 2154 1961 2206
rect 3209 2154 3261 2206
rect 3474 2154 3526 2206
rect 3604 2154 3656 2206
rect 3734 2154 3786 2206
rect 4254 2154 4306 2206
rect 4384 2154 4436 2206
rect 4504 2154 4556 2206
rect 184 1964 236 2016
rect 184 1874 236 1926
rect 444 1964 496 2016
rect 444 1874 496 1926
rect 704 1964 756 2016
rect 704 1874 756 1926
rect 964 1964 1016 2016
rect 964 1874 1016 1926
rect 1224 1964 1276 2016
rect 1224 1874 1276 1926
rect 1484 1964 1536 2016
rect 1484 1874 1536 1926
rect 1744 1964 1796 2016
rect 1744 1874 1796 1926
rect 2004 1964 2056 2016
rect 2004 1874 2056 1926
rect 2264 1964 2316 2016
rect 2264 1874 2316 1926
rect 2524 1964 2576 2016
rect 2524 1874 2576 1926
rect 2784 1964 2836 2016
rect 2784 1874 2836 1926
rect 3044 1964 3096 2016
rect 3044 1874 3096 1926
rect 3304 1964 3356 2016
rect 3304 1874 3356 1926
rect 3564 1964 3616 2016
rect 3564 1874 3616 1926
rect 3824 1964 3876 2016
rect 3824 1874 3876 1926
rect 4084 1964 4136 2016
rect 4084 1874 4136 1926
rect 4344 1964 4396 2016
rect 4344 1874 4396 1926
rect 4604 1964 4656 2016
rect 4604 1874 4656 1926
rect 4864 1964 4916 2016
rect 4864 1874 4916 1926
rect 5124 1964 5176 2016
rect 5124 1874 5176 1926
rect -171 94 -119 146
rect -41 94 11 146
rect 89 94 141 146
rect 349 94 401 146
rect 609 94 661 146
rect 609 -176 661 -124
rect 869 94 921 146
rect 869 -176 921 -124
rect 1129 94 1181 146
rect 1389 94 1441 146
rect 1389 -176 1441 -124
rect 1649 94 1701 146
rect 1649 -176 1701 -124
rect 1909 94 1961 146
rect 1909 -176 1961 -124
rect 2169 94 2221 146
rect 2429 94 2481 146
rect 2689 94 2741 146
rect 2949 94 3001 146
rect 3209 94 3261 146
rect 3209 -176 3261 -124
rect 3469 94 3521 146
rect 3469 -176 3521 -124
rect 3729 94 3781 146
rect 3729 -176 3781 -124
rect 3989 94 4041 146
rect 4249 94 4301 146
rect 4249 -176 4301 -124
rect 4509 94 4561 146
rect 4509 -176 4561 -124
rect 4769 94 4821 146
rect 5029 94 5081 146
rect 5254 94 5306 146
rect 5334 94 5386 146
rect 5394 -86 5446 -34
rect 5474 -86 5526 -34
rect -171 -2236 -119 -2184
rect -81 -2236 -29 -2184
rect 89 -2236 141 -2184
rect 349 -2236 401 -2184
rect 609 -2236 661 -2184
rect 869 -2236 921 -2184
rect 1129 -2236 1181 -2184
rect 1389 -2236 1441 -2184
rect 1649 -2236 1701 -2184
rect 1909 -2236 1961 -2184
rect 2169 -2236 2221 -2184
rect 2429 -2236 2481 -2184
rect 2689 -2236 2741 -2184
rect 2949 -2236 3001 -2184
rect 3209 -2236 3261 -2184
rect 3469 -2236 3521 -2184
rect 3729 -2236 3781 -2184
rect 3989 -2236 4041 -2184
rect 4249 -2236 4301 -2184
rect 4509 -2236 4561 -2184
rect 4769 -2236 4821 -2184
rect 5029 -2236 5081 -2184
rect 5144 -2236 5196 -2184
rect 5274 -2236 5326 -2184
rect -286 -2416 -234 -2364
rect -206 -2416 -154 -2364
rect 5574 -2236 5626 -2184
rect 5574 -2316 5626 -2264
rect 5664 -6 5716 46
rect 5664 -86 5716 -34
rect 5394 -2416 5446 -2364
rect 5474 -2416 5526 -2364
rect 5574 -2736 5626 -2684
rect 5654 -2736 5706 -2684
rect -466 -2826 -414 -2774
rect -386 -2826 -334 -2774
<< metal2 >>
rect -390 2808 -220 2820
rect -390 2752 -378 2808
rect -322 2752 -288 2808
rect -232 2800 -220 2808
rect 5570 2808 5740 2820
rect 5570 2800 5582 2808
rect -232 2752 5582 2800
rect 5638 2752 5672 2808
rect 5728 2752 5740 2808
rect -390 2740 5740 2752
rect -390 2706 6130 2710
rect -390 2654 -376 2706
rect -324 2698 6130 2706
rect -324 2654 5352 2698
rect -390 2650 5352 2654
rect 5340 2642 5352 2650
rect 5408 2642 5442 2698
rect 5498 2650 6130 2698
rect 5498 2642 5510 2650
rect 5340 2630 5510 2642
rect 6030 2618 6130 2650
rect 6030 2562 6052 2618
rect 6108 2562 6130 2618
rect 6030 2540 6130 2562
rect -530 2378 1940 2390
rect -530 2322 -518 2378
rect -462 2330 1940 2378
rect -462 2322 -450 2330
rect -530 2288 -450 2322
rect -530 2232 -518 2288
rect -462 2232 -450 2288
rect -530 2220 -450 2232
rect -390 2286 -330 2300
rect -390 2234 -386 2286
rect -334 2234 -330 2286
rect -300 2296 1730 2300
rect -300 2244 -286 2296
rect -234 2244 -206 2296
rect -154 2244 1730 2296
rect -300 2240 1730 2244
rect -390 2210 -330 2234
rect -390 2206 940 2210
rect -390 2154 -386 2206
rect -334 2154 604 2206
rect 656 2154 704 2206
rect 756 2154 804 2206
rect 856 2154 940 2206
rect -390 2150 940 2154
rect 1370 2206 1730 2240
rect 1370 2154 1394 2206
rect 1446 2154 1514 2206
rect 1566 2154 1634 2206
rect 1686 2154 1730 2206
rect 1370 2150 1730 2154
rect 1890 2210 1940 2330
rect 3220 2330 5740 2390
rect 3220 2210 3280 2330
rect 1890 2206 1980 2210
rect 1890 2154 1909 2206
rect 1961 2154 1980 2206
rect 1890 2150 1980 2154
rect 3190 2206 3280 2210
rect 3190 2154 3209 2206
rect 3261 2154 3280 2206
rect 3190 2150 3280 2154
rect 3450 2296 5630 2300
rect 3450 2244 5484 2296
rect 5536 2244 5564 2296
rect 5616 2244 5630 2296
rect 3450 2240 5630 2244
rect 3450 2206 3800 2240
rect 3450 2154 3474 2206
rect 3526 2154 3604 2206
rect 3656 2154 3734 2206
rect 3786 2154 3800 2206
rect 3450 2150 3800 2154
rect 4230 2206 5650 2210
rect 4230 2154 4254 2206
rect 4306 2154 4384 2206
rect 4436 2154 4504 2206
rect 4556 2198 5650 2206
rect 4556 2154 5582 2198
rect 4230 2150 5582 2154
rect -390 2140 -330 2150
rect 5570 2142 5582 2150
rect 5638 2142 5650 2198
rect 5570 2108 5650 2142
rect 5570 2052 5582 2108
rect 5638 2052 5650 2108
rect 5570 2040 5650 2052
rect 170 2018 250 2030
rect 170 1962 182 2018
rect 238 1962 250 2018
rect 170 1928 250 1962
rect 170 1872 182 1928
rect 238 1872 250 1928
rect 170 1860 250 1872
rect 430 2018 510 2030
rect 430 1962 442 2018
rect 498 1962 510 2018
rect 430 1928 510 1962
rect 430 1872 442 1928
rect 498 1872 510 1928
rect 430 1860 510 1872
rect 690 2018 770 2030
rect 690 1962 702 2018
rect 758 1962 770 2018
rect 690 1928 770 1962
rect 690 1872 702 1928
rect 758 1872 770 1928
rect 690 1860 770 1872
rect 950 2018 1030 2030
rect 950 1962 962 2018
rect 1018 1962 1030 2018
rect 950 1928 1030 1962
rect 950 1872 962 1928
rect 1018 1872 1030 1928
rect 950 1860 1030 1872
rect 1210 2018 1290 2030
rect 1210 1962 1222 2018
rect 1278 1962 1290 2018
rect 1210 1928 1290 1962
rect 1210 1872 1222 1928
rect 1278 1872 1290 1928
rect 1210 1860 1290 1872
rect 1470 2018 1550 2030
rect 1470 1962 1482 2018
rect 1538 1962 1550 2018
rect 1470 1928 1550 1962
rect 1470 1872 1482 1928
rect 1538 1872 1550 1928
rect 1470 1860 1550 1872
rect 1730 2018 1810 2030
rect 1730 1962 1742 2018
rect 1798 1962 1810 2018
rect 1730 1928 1810 1962
rect 1730 1872 1742 1928
rect 1798 1872 1810 1928
rect 1730 1860 1810 1872
rect 1990 2018 2070 2030
rect 1990 1962 2002 2018
rect 2058 1962 2070 2018
rect 1990 1928 2070 1962
rect 1990 1872 2002 1928
rect 2058 1872 2070 1928
rect 1990 1860 2070 1872
rect 2250 2018 2330 2030
rect 2250 1962 2262 2018
rect 2318 1962 2330 2018
rect 2250 1928 2330 1962
rect 2250 1872 2262 1928
rect 2318 1872 2330 1928
rect 2250 1860 2330 1872
rect 2510 2018 2590 2030
rect 2510 1962 2522 2018
rect 2578 1962 2590 2018
rect 2510 1928 2590 1962
rect 2510 1872 2522 1928
rect 2578 1872 2590 1928
rect 2510 1860 2590 1872
rect 2770 2018 2850 2030
rect 2770 1962 2782 2018
rect 2838 1962 2850 2018
rect 2770 1928 2850 1962
rect 2770 1872 2782 1928
rect 2838 1872 2850 1928
rect 2770 1860 2850 1872
rect 3030 2018 3110 2030
rect 3030 1962 3042 2018
rect 3098 1962 3110 2018
rect 3030 1928 3110 1962
rect 3030 1872 3042 1928
rect 3098 1872 3110 1928
rect 3030 1860 3110 1872
rect 3290 2018 3370 2030
rect 3290 1962 3302 2018
rect 3358 1962 3370 2018
rect 3290 1928 3370 1962
rect 3290 1872 3302 1928
rect 3358 1872 3370 1928
rect 3290 1860 3370 1872
rect 3550 2018 3630 2030
rect 3550 1962 3562 2018
rect 3618 1962 3630 2018
rect 3550 1928 3630 1962
rect 3550 1872 3562 1928
rect 3618 1872 3630 1928
rect 3550 1860 3630 1872
rect 3810 2018 3890 2030
rect 3810 1962 3822 2018
rect 3878 1962 3890 2018
rect 3810 1928 3890 1962
rect 3810 1872 3822 1928
rect 3878 1872 3890 1928
rect 3810 1860 3890 1872
rect 4070 2018 4150 2030
rect 4070 1962 4082 2018
rect 4138 1962 4150 2018
rect 4070 1928 4150 1962
rect 4070 1872 4082 1928
rect 4138 1872 4150 1928
rect 4070 1860 4150 1872
rect 4330 2018 4410 2030
rect 4330 1962 4342 2018
rect 4398 1962 4410 2018
rect 4330 1928 4410 1962
rect 4330 1872 4342 1928
rect 4398 1872 4410 1928
rect 4330 1860 4410 1872
rect 4590 2018 4670 2030
rect 4590 1962 4602 2018
rect 4658 1962 4670 2018
rect 4590 1928 4670 1962
rect 4590 1872 4602 1928
rect 4658 1872 4670 1928
rect 4590 1860 4670 1872
rect 4850 2018 4930 2030
rect 4850 1962 4862 2018
rect 4918 1962 4930 2018
rect 4850 1928 4930 1962
rect 4850 1872 4862 1928
rect 4918 1872 4930 1928
rect 4850 1860 4930 1872
rect 5110 2018 5190 2030
rect 5110 1962 5122 2018
rect 5178 1962 5190 2018
rect 5110 1928 5190 1962
rect 5110 1872 5122 1928
rect 5178 1872 5190 1928
rect 5110 1860 5190 1872
rect 5680 1980 5740 2330
rect 5680 1968 5760 1980
rect 5680 1912 5692 1968
rect 5748 1912 5760 1968
rect 5680 1878 5760 1912
rect 5680 1822 5692 1878
rect 5748 1822 5760 1878
rect 5680 1810 5760 1822
rect -190 146 5400 150
rect -190 94 -171 146
rect -119 94 -41 146
rect 11 94 89 146
rect 141 94 349 146
rect 401 94 609 146
rect 661 94 869 146
rect 921 94 1129 146
rect 1181 94 1389 146
rect 1441 94 1649 146
rect 1701 94 1909 146
rect 1961 94 2169 146
rect 2221 94 2429 146
rect 2481 94 2689 146
rect 2741 94 2949 146
rect 3001 94 3209 146
rect 3261 94 3469 146
rect 3521 94 3729 146
rect 3781 94 3989 146
rect 4041 94 4249 146
rect 4301 94 4509 146
rect 4561 94 4769 146
rect 4821 94 5029 146
rect 5081 94 5254 146
rect 5306 94 5334 146
rect 5386 94 5400 146
rect -190 90 5400 94
rect -480 46 1950 60
rect -480 -6 -476 46
rect -424 0 1950 46
rect -424 -6 -420 0
rect -480 -34 -420 -6
rect -480 -86 -476 -34
rect -424 -86 -420 -34
rect -480 -100 -420 -86
rect -390 -44 1720 -30
rect -390 -96 -386 -44
rect -334 -90 1720 -44
rect -334 -96 -330 -90
rect -390 -124 -330 -96
rect -390 -176 -386 -124
rect -334 -176 -330 -124
rect -390 -190 -330 -176
rect -300 -124 940 -120
rect -300 -132 609 -124
rect -300 -188 -288 -132
rect -232 -176 609 -132
rect 661 -176 869 -124
rect 921 -176 940 -124
rect -232 -180 940 -176
rect 1370 -124 1720 -90
rect 1370 -176 1389 -124
rect 1441 -176 1649 -124
rect 1701 -176 1720 -124
rect 1370 -180 1720 -176
rect 1890 -120 1950 0
rect 3190 46 5720 60
rect 3190 0 5664 46
rect 1890 -124 1980 -120
rect 1890 -176 1909 -124
rect 1961 -176 1980 -124
rect 1890 -180 1980 -176
rect 3190 -124 3280 0
rect 5660 -6 5664 0
rect 5716 -6 5720 46
rect 3190 -176 3209 -124
rect 3261 -176 3280 -124
rect 3190 -180 3280 -176
rect 3450 -34 5540 -30
rect 3450 -86 5394 -34
rect 5446 -86 5474 -34
rect 5526 -86 5540 -34
rect 3450 -90 5540 -86
rect 5660 -34 5720 -6
rect 5660 -86 5664 -34
rect 5716 -86 5720 -34
rect 3450 -124 3810 -90
rect 5660 -100 5720 -86
rect 3450 -176 3469 -124
rect 3521 -176 3729 -124
rect 3781 -176 3810 -124
rect 3450 -180 3810 -176
rect 4230 -124 5540 -120
rect 4230 -176 4249 -124
rect 4301 -176 4509 -124
rect 4561 -132 5540 -124
rect 4561 -176 5382 -132
rect 4230 -180 5382 -176
rect -232 -188 -220 -180
rect -300 -200 -220 -188
rect 5370 -188 5382 -180
rect 5438 -188 5472 -132
rect 5528 -188 5540 -132
rect 5370 -200 5540 -188
rect -390 -2184 -330 -2170
rect -390 -2236 -386 -2184
rect -334 -2236 -330 -2184
rect -390 -2264 -330 -2236
rect -190 -2184 5360 -2180
rect -190 -2236 -171 -2184
rect -119 -2236 -81 -2184
rect -29 -2236 89 -2184
rect 141 -2236 349 -2184
rect 401 -2236 609 -2184
rect 661 -2236 869 -2184
rect 921 -2236 1129 -2184
rect 1181 -2236 1389 -2184
rect 1441 -2236 1649 -2184
rect 1701 -2236 1909 -2184
rect 1961 -2236 2169 -2184
rect 2221 -2236 2429 -2184
rect 2481 -2236 2689 -2184
rect 2741 -2236 2949 -2184
rect 3001 -2236 3209 -2184
rect 3261 -2236 3469 -2184
rect 3521 -2236 3729 -2184
rect 3781 -2236 3989 -2184
rect 4041 -2236 4249 -2184
rect 4301 -2236 4509 -2184
rect 4561 -2236 4769 -2184
rect 4821 -2236 5029 -2184
rect 5081 -2236 5144 -2184
rect 5196 -2236 5274 -2184
rect 5326 -2236 5360 -2184
rect -190 -2240 5360 -2236
rect 5570 -2184 5630 -2170
rect 5570 -2236 5574 -2184
rect 5626 -2236 5630 -2184
rect -390 -2316 -386 -2264
rect -334 -2270 -330 -2264
rect 5570 -2264 5630 -2236
rect 5570 -2270 5574 -2264
rect -334 -2316 5574 -2270
rect 5626 -2270 5630 -2264
rect 6030 -2182 6130 -2160
rect 6030 -2238 6052 -2182
rect 6108 -2238 6130 -2182
rect 6030 -2270 6130 -2238
rect 5626 -2316 6130 -2270
rect -390 -2330 6130 -2316
rect -300 -2364 6130 -2360
rect -300 -2416 -286 -2364
rect -234 -2416 -206 -2364
rect -154 -2416 5394 -2364
rect 5446 -2416 5474 -2364
rect 5526 -2382 6130 -2364
rect 5526 -2416 6052 -2382
rect -300 -2420 6052 -2416
rect 6030 -2438 6052 -2420
rect 6108 -2438 6130 -2382
rect 6030 -2460 6130 -2438
rect -510 -2582 -430 -2570
rect -510 -2638 -498 -2582
rect -442 -2638 -430 -2582
rect 6030 -2602 6130 -2580
rect 6030 -2630 6052 -2602
rect -510 -2672 -430 -2638
rect -510 -2728 -498 -2672
rect -442 -2680 -430 -2672
rect 5660 -2658 6052 -2630
rect 6108 -2658 6130 -2602
rect 5660 -2680 6130 -2658
rect -442 -2684 5720 -2680
rect -442 -2728 5574 -2684
rect -510 -2736 5574 -2728
rect 5626 -2736 5654 -2684
rect 5706 -2736 5720 -2684
rect -510 -2740 5720 -2736
rect -480 -2774 5760 -2770
rect -480 -2826 -466 -2774
rect -414 -2826 -386 -2774
rect -334 -2782 5760 -2774
rect -334 -2826 5602 -2782
rect -480 -2830 5602 -2826
rect 5590 -2838 5602 -2830
rect 5658 -2838 5692 -2782
rect 5748 -2838 5760 -2782
rect 5590 -2850 5760 -2838
<< via2 >>
rect -378 2752 -322 2808
rect -288 2752 -232 2808
rect 5582 2752 5638 2808
rect 5672 2752 5728 2808
rect 5352 2642 5408 2698
rect 5442 2642 5498 2698
rect 6052 2562 6108 2618
rect -518 2322 -462 2378
rect -518 2232 -462 2288
rect 5582 2142 5638 2198
rect 5582 2052 5638 2108
rect 182 2016 238 2018
rect 182 1964 184 2016
rect 184 1964 236 2016
rect 236 1964 238 2016
rect 182 1962 238 1964
rect 182 1926 238 1928
rect 182 1874 184 1926
rect 184 1874 236 1926
rect 236 1874 238 1926
rect 182 1872 238 1874
rect 442 2016 498 2018
rect 442 1964 444 2016
rect 444 1964 496 2016
rect 496 1964 498 2016
rect 442 1962 498 1964
rect 442 1926 498 1928
rect 442 1874 444 1926
rect 444 1874 496 1926
rect 496 1874 498 1926
rect 442 1872 498 1874
rect 702 2016 758 2018
rect 702 1964 704 2016
rect 704 1964 756 2016
rect 756 1964 758 2016
rect 702 1962 758 1964
rect 702 1926 758 1928
rect 702 1874 704 1926
rect 704 1874 756 1926
rect 756 1874 758 1926
rect 702 1872 758 1874
rect 962 2016 1018 2018
rect 962 1964 964 2016
rect 964 1964 1016 2016
rect 1016 1964 1018 2016
rect 962 1962 1018 1964
rect 962 1926 1018 1928
rect 962 1874 964 1926
rect 964 1874 1016 1926
rect 1016 1874 1018 1926
rect 962 1872 1018 1874
rect 1222 2016 1278 2018
rect 1222 1964 1224 2016
rect 1224 1964 1276 2016
rect 1276 1964 1278 2016
rect 1222 1962 1278 1964
rect 1222 1926 1278 1928
rect 1222 1874 1224 1926
rect 1224 1874 1276 1926
rect 1276 1874 1278 1926
rect 1222 1872 1278 1874
rect 1482 2016 1538 2018
rect 1482 1964 1484 2016
rect 1484 1964 1536 2016
rect 1536 1964 1538 2016
rect 1482 1962 1538 1964
rect 1482 1926 1538 1928
rect 1482 1874 1484 1926
rect 1484 1874 1536 1926
rect 1536 1874 1538 1926
rect 1482 1872 1538 1874
rect 1742 2016 1798 2018
rect 1742 1964 1744 2016
rect 1744 1964 1796 2016
rect 1796 1964 1798 2016
rect 1742 1962 1798 1964
rect 1742 1926 1798 1928
rect 1742 1874 1744 1926
rect 1744 1874 1796 1926
rect 1796 1874 1798 1926
rect 1742 1872 1798 1874
rect 2002 2016 2058 2018
rect 2002 1964 2004 2016
rect 2004 1964 2056 2016
rect 2056 1964 2058 2016
rect 2002 1962 2058 1964
rect 2002 1926 2058 1928
rect 2002 1874 2004 1926
rect 2004 1874 2056 1926
rect 2056 1874 2058 1926
rect 2002 1872 2058 1874
rect 2262 2016 2318 2018
rect 2262 1964 2264 2016
rect 2264 1964 2316 2016
rect 2316 1964 2318 2016
rect 2262 1962 2318 1964
rect 2262 1926 2318 1928
rect 2262 1874 2264 1926
rect 2264 1874 2316 1926
rect 2316 1874 2318 1926
rect 2262 1872 2318 1874
rect 2522 2016 2578 2018
rect 2522 1964 2524 2016
rect 2524 1964 2576 2016
rect 2576 1964 2578 2016
rect 2522 1962 2578 1964
rect 2522 1926 2578 1928
rect 2522 1874 2524 1926
rect 2524 1874 2576 1926
rect 2576 1874 2578 1926
rect 2522 1872 2578 1874
rect 2782 2016 2838 2018
rect 2782 1964 2784 2016
rect 2784 1964 2836 2016
rect 2836 1964 2838 2016
rect 2782 1962 2838 1964
rect 2782 1926 2838 1928
rect 2782 1874 2784 1926
rect 2784 1874 2836 1926
rect 2836 1874 2838 1926
rect 2782 1872 2838 1874
rect 3042 2016 3098 2018
rect 3042 1964 3044 2016
rect 3044 1964 3096 2016
rect 3096 1964 3098 2016
rect 3042 1962 3098 1964
rect 3042 1926 3098 1928
rect 3042 1874 3044 1926
rect 3044 1874 3096 1926
rect 3096 1874 3098 1926
rect 3042 1872 3098 1874
rect 3302 2016 3358 2018
rect 3302 1964 3304 2016
rect 3304 1964 3356 2016
rect 3356 1964 3358 2016
rect 3302 1962 3358 1964
rect 3302 1926 3358 1928
rect 3302 1874 3304 1926
rect 3304 1874 3356 1926
rect 3356 1874 3358 1926
rect 3302 1872 3358 1874
rect 3562 2016 3618 2018
rect 3562 1964 3564 2016
rect 3564 1964 3616 2016
rect 3616 1964 3618 2016
rect 3562 1962 3618 1964
rect 3562 1926 3618 1928
rect 3562 1874 3564 1926
rect 3564 1874 3616 1926
rect 3616 1874 3618 1926
rect 3562 1872 3618 1874
rect 3822 2016 3878 2018
rect 3822 1964 3824 2016
rect 3824 1964 3876 2016
rect 3876 1964 3878 2016
rect 3822 1962 3878 1964
rect 3822 1926 3878 1928
rect 3822 1874 3824 1926
rect 3824 1874 3876 1926
rect 3876 1874 3878 1926
rect 3822 1872 3878 1874
rect 4082 2016 4138 2018
rect 4082 1964 4084 2016
rect 4084 1964 4136 2016
rect 4136 1964 4138 2016
rect 4082 1962 4138 1964
rect 4082 1926 4138 1928
rect 4082 1874 4084 1926
rect 4084 1874 4136 1926
rect 4136 1874 4138 1926
rect 4082 1872 4138 1874
rect 4342 2016 4398 2018
rect 4342 1964 4344 2016
rect 4344 1964 4396 2016
rect 4396 1964 4398 2016
rect 4342 1962 4398 1964
rect 4342 1926 4398 1928
rect 4342 1874 4344 1926
rect 4344 1874 4396 1926
rect 4396 1874 4398 1926
rect 4342 1872 4398 1874
rect 4602 2016 4658 2018
rect 4602 1964 4604 2016
rect 4604 1964 4656 2016
rect 4656 1964 4658 2016
rect 4602 1962 4658 1964
rect 4602 1926 4658 1928
rect 4602 1874 4604 1926
rect 4604 1874 4656 1926
rect 4656 1874 4658 1926
rect 4602 1872 4658 1874
rect 4862 2016 4918 2018
rect 4862 1964 4864 2016
rect 4864 1964 4916 2016
rect 4916 1964 4918 2016
rect 4862 1962 4918 1964
rect 4862 1926 4918 1928
rect 4862 1874 4864 1926
rect 4864 1874 4916 1926
rect 4916 1874 4918 1926
rect 4862 1872 4918 1874
rect 5122 2016 5178 2018
rect 5122 1964 5124 2016
rect 5124 1964 5176 2016
rect 5176 1964 5178 2016
rect 5122 1962 5178 1964
rect 5122 1926 5178 1928
rect 5122 1874 5124 1926
rect 5124 1874 5176 1926
rect 5176 1874 5178 1926
rect 5122 1872 5178 1874
rect 5692 1912 5748 1968
rect 5692 1822 5748 1878
rect -288 -188 -232 -132
rect 5382 -188 5438 -132
rect 5472 -188 5528 -132
rect 6052 -2238 6108 -2182
rect 6052 -2438 6108 -2382
rect -498 -2638 -442 -2582
rect -498 -2728 -442 -2672
rect 6052 -2658 6108 -2602
rect 5602 -2838 5658 -2782
rect 5692 -2838 5748 -2782
<< metal3 >>
rect 170 2912 270 2930
rect 170 2848 188 2912
rect 252 2848 270 2912
rect 170 2830 270 2848
rect 430 2912 530 2930
rect 430 2848 448 2912
rect 512 2848 530 2912
rect 430 2830 530 2848
rect 690 2912 790 2930
rect 690 2848 708 2912
rect 772 2848 790 2912
rect 690 2830 790 2848
rect 950 2912 1050 2930
rect 950 2848 968 2912
rect 1032 2848 1050 2912
rect 950 2830 1050 2848
rect 1210 2912 1310 2930
rect 1210 2848 1228 2912
rect 1292 2848 1310 2912
rect 1210 2830 1310 2848
rect 1470 2912 1570 2930
rect 1470 2848 1488 2912
rect 1552 2848 1570 2912
rect 1470 2830 1570 2848
rect 1730 2912 1830 2930
rect 1730 2848 1748 2912
rect 1812 2848 1830 2912
rect 1730 2830 1830 2848
rect 1990 2912 2090 2930
rect 1990 2848 2008 2912
rect 2072 2848 2090 2912
rect 1990 2830 2090 2848
rect 2250 2912 2350 2930
rect 2250 2848 2268 2912
rect 2332 2848 2350 2912
rect 2250 2830 2350 2848
rect 2510 2912 2610 2930
rect 2510 2848 2528 2912
rect 2592 2848 2610 2912
rect 2510 2830 2610 2848
rect 2770 2912 2870 2930
rect 2770 2848 2788 2912
rect 2852 2848 2870 2912
rect 2770 2830 2870 2848
rect 3030 2912 3130 2930
rect 3030 2848 3048 2912
rect 3112 2848 3130 2912
rect 3030 2830 3130 2848
rect 3290 2912 3390 2930
rect 3290 2848 3308 2912
rect 3372 2848 3390 2912
rect 3290 2830 3390 2848
rect 3550 2912 3650 2930
rect 3550 2848 3568 2912
rect 3632 2848 3650 2912
rect 3550 2830 3650 2848
rect 3810 2912 3910 2930
rect 3810 2848 3828 2912
rect 3892 2848 3910 2912
rect 3810 2830 3910 2848
rect 4070 2912 4170 2930
rect 4070 2848 4088 2912
rect 4152 2848 4170 2912
rect 4070 2830 4170 2848
rect 4330 2912 4430 2930
rect 4330 2848 4348 2912
rect 4412 2848 4430 2912
rect 4330 2830 4430 2848
rect 4590 2912 4690 2930
rect 4590 2848 4608 2912
rect 4672 2848 4690 2912
rect 4590 2830 4690 2848
rect 4850 2912 4950 2930
rect 4850 2848 4868 2912
rect 4932 2848 4950 2912
rect 4850 2830 4950 2848
rect 5110 2912 5210 2930
rect 5110 2848 5128 2912
rect 5192 2848 5210 2912
rect 5110 2830 5210 2848
rect -390 2808 -220 2820
rect -390 2752 -378 2808
rect -322 2752 -288 2808
rect -232 2752 -220 2808
rect -390 2740 -220 2752
rect -530 2378 -450 2390
rect -530 2322 -518 2378
rect -462 2322 -450 2378
rect -530 2288 -450 2322
rect -530 2232 -518 2288
rect -462 2232 -450 2288
rect -530 2220 -450 2232
rect -510 -2570 -450 2220
rect -390 -120 -330 2740
rect 190 2030 250 2830
rect 450 2030 510 2830
rect 710 2030 770 2830
rect 970 2030 1030 2830
rect 1230 2030 1290 2830
rect 1490 2030 1550 2830
rect 1750 2030 1810 2830
rect 2010 2030 2070 2830
rect 2270 2030 2330 2830
rect 2530 2030 2590 2830
rect 2790 2030 2850 2830
rect 3050 2030 3110 2830
rect 3310 2030 3370 2830
rect 3570 2030 3630 2830
rect 3830 2030 3890 2830
rect 4090 2030 4150 2830
rect 4350 2030 4410 2830
rect 4610 2030 4670 2830
rect 4870 2030 4930 2830
rect 5130 2030 5190 2830
rect 6030 2820 6130 2840
rect 5570 2808 6130 2820
rect 5570 2752 5582 2808
rect 5638 2752 5672 2808
rect 5728 2752 6130 2808
rect 5570 2740 6130 2752
rect 5340 2698 5510 2710
rect 5340 2642 5352 2698
rect 5408 2642 5442 2698
rect 5498 2642 5510 2698
rect 5340 2630 5510 2642
rect 170 2018 250 2030
rect 170 1962 182 2018
rect 238 1962 250 2018
rect 170 1928 250 1962
rect 170 1872 182 1928
rect 238 1872 250 1928
rect 170 1860 250 1872
rect 430 2018 510 2030
rect 430 1962 442 2018
rect 498 1962 510 2018
rect 430 1928 510 1962
rect 430 1872 442 1928
rect 498 1872 510 1928
rect 430 1860 510 1872
rect 690 2018 770 2030
rect 690 1962 702 2018
rect 758 1962 770 2018
rect 690 1928 770 1962
rect 690 1872 702 1928
rect 758 1872 770 1928
rect 690 1860 770 1872
rect 950 2018 1030 2030
rect 950 1962 962 2018
rect 1018 1962 1030 2018
rect 950 1928 1030 1962
rect 950 1872 962 1928
rect 1018 1872 1030 1928
rect 950 1860 1030 1872
rect 1210 2018 1290 2030
rect 1210 1962 1222 2018
rect 1278 1962 1290 2018
rect 1210 1928 1290 1962
rect 1210 1872 1222 1928
rect 1278 1872 1290 1928
rect 1210 1860 1290 1872
rect 1470 2018 1550 2030
rect 1470 1962 1482 2018
rect 1538 1962 1550 2018
rect 1470 1928 1550 1962
rect 1470 1872 1482 1928
rect 1538 1872 1550 1928
rect 1470 1860 1550 1872
rect 1730 2018 1810 2030
rect 1730 1962 1742 2018
rect 1798 1962 1810 2018
rect 1730 1928 1810 1962
rect 1730 1872 1742 1928
rect 1798 1872 1810 1928
rect 1730 1860 1810 1872
rect 1990 2018 2070 2030
rect 1990 1962 2002 2018
rect 2058 1962 2070 2018
rect 1990 1928 2070 1962
rect 1990 1872 2002 1928
rect 2058 1872 2070 1928
rect 1990 1860 2070 1872
rect 2250 2018 2330 2030
rect 2250 1962 2262 2018
rect 2318 1962 2330 2018
rect 2250 1928 2330 1962
rect 2250 1872 2262 1928
rect 2318 1872 2330 1928
rect 2250 1860 2330 1872
rect 2510 2018 2590 2030
rect 2510 1962 2522 2018
rect 2578 1962 2590 2018
rect 2510 1928 2590 1962
rect 2510 1872 2522 1928
rect 2578 1872 2590 1928
rect 2510 1860 2590 1872
rect 2770 2018 2850 2030
rect 2770 1962 2782 2018
rect 2838 1962 2850 2018
rect 2770 1928 2850 1962
rect 2770 1872 2782 1928
rect 2838 1872 2850 1928
rect 2770 1860 2850 1872
rect 3030 2018 3110 2030
rect 3030 1962 3042 2018
rect 3098 1962 3110 2018
rect 3030 1928 3110 1962
rect 3030 1872 3042 1928
rect 3098 1872 3110 1928
rect 3030 1860 3110 1872
rect 3290 2018 3370 2030
rect 3290 1962 3302 2018
rect 3358 1962 3370 2018
rect 3290 1928 3370 1962
rect 3290 1872 3302 1928
rect 3358 1872 3370 1928
rect 3290 1860 3370 1872
rect 3550 2018 3630 2030
rect 3550 1962 3562 2018
rect 3618 1962 3630 2018
rect 3550 1928 3630 1962
rect 3550 1872 3562 1928
rect 3618 1872 3630 1928
rect 3550 1860 3630 1872
rect 3810 2018 3890 2030
rect 3810 1962 3822 2018
rect 3878 1962 3890 2018
rect 3810 1928 3890 1962
rect 3810 1872 3822 1928
rect 3878 1872 3890 1928
rect 3810 1860 3890 1872
rect 4070 2018 4150 2030
rect 4070 1962 4082 2018
rect 4138 1962 4150 2018
rect 4070 1928 4150 1962
rect 4070 1872 4082 1928
rect 4138 1872 4150 1928
rect 4070 1860 4150 1872
rect 4330 2018 4410 2030
rect 4330 1962 4342 2018
rect 4398 1962 4410 2018
rect 4330 1928 4410 1962
rect 4330 1872 4342 1928
rect 4398 1872 4410 1928
rect 4330 1860 4410 1872
rect 4590 2018 4670 2030
rect 4590 1962 4602 2018
rect 4658 1962 4670 2018
rect 4590 1928 4670 1962
rect 4590 1872 4602 1928
rect 4658 1872 4670 1928
rect 4590 1860 4670 1872
rect 4850 2018 4930 2030
rect 4850 1962 4862 2018
rect 4918 1962 4930 2018
rect 4850 1928 4930 1962
rect 4850 1872 4862 1928
rect 4918 1872 4930 1928
rect 4850 1860 4930 1872
rect 5110 2018 5190 2030
rect 5110 1962 5122 2018
rect 5178 1962 5190 2018
rect 5110 1928 5190 1962
rect 5110 1872 5122 1928
rect 5178 1872 5190 1928
rect 5110 1860 5190 1872
rect 5450 -120 5510 2630
rect 5570 2210 5630 2740
rect 6030 2618 6130 2640
rect 6030 2562 6052 2618
rect 6108 2562 6130 2618
rect 6030 2540 6130 2562
rect 5570 2198 5650 2210
rect 5570 2142 5582 2198
rect 5638 2142 5650 2198
rect 5570 2108 5650 2142
rect 5570 2052 5582 2108
rect 5638 2052 5650 2108
rect 5570 2040 5650 2052
rect 5680 1968 5760 1980
rect 5680 1912 5692 1968
rect 5748 1912 5760 1968
rect 5680 1878 5760 1912
rect 5680 1822 5692 1878
rect 5748 1822 5760 1878
rect -390 -132 -220 -120
rect -390 -180 -288 -132
rect -300 -188 -288 -180
rect -232 -188 -220 -132
rect -300 -200 -220 -188
rect 5370 -132 5540 -120
rect 5370 -188 5382 -132
rect 5438 -188 5472 -132
rect 5528 -188 5540 -132
rect 5370 -200 5540 -188
rect -510 -2582 -430 -2570
rect -510 -2638 -498 -2582
rect -442 -2638 -430 -2582
rect -510 -2672 -430 -2638
rect -510 -2728 -498 -2672
rect -442 -2728 -430 -2672
rect -510 -2740 -430 -2728
rect 5680 -2770 5760 1822
rect 6030 -2182 6130 -2160
rect 6030 -2238 6052 -2182
rect 6108 -2238 6130 -2182
rect 6030 -2260 6130 -2238
rect 6040 -2382 6120 -2370
rect 6040 -2438 6052 -2382
rect 6108 -2438 6120 -2382
rect 6040 -2450 6120 -2438
rect 6030 -2602 6130 -2580
rect 6030 -2658 6052 -2602
rect 6108 -2658 6130 -2602
rect 6030 -2680 6130 -2658
rect 5590 -2782 6130 -2770
rect 5590 -2838 5602 -2782
rect 5658 -2838 5692 -2782
rect 5748 -2838 6130 -2782
rect 5590 -2850 6130 -2838
rect 6030 -2870 6130 -2850
<< via3 >>
rect 188 2848 252 2912
rect 448 2848 512 2912
rect 708 2848 772 2912
rect 968 2848 1032 2912
rect 1228 2848 1292 2912
rect 1488 2848 1552 2912
rect 1748 2848 1812 2912
rect 2008 2848 2072 2912
rect 2268 2848 2332 2912
rect 2528 2848 2592 2912
rect 2788 2848 2852 2912
rect 3048 2848 3112 2912
rect 3308 2848 3372 2912
rect 3568 2848 3632 2912
rect 3828 2848 3892 2912
rect 4088 2848 4152 2912
rect 4348 2848 4412 2912
rect 4608 2848 4672 2912
rect 4868 2848 4932 2912
rect 5128 2848 5192 2912
<< metal4 >>
rect -770 2912 5470 2930
rect -770 2848 188 2912
rect 252 2848 448 2912
rect 512 2848 708 2912
rect 772 2848 968 2912
rect 1032 2848 1228 2912
rect 1292 2848 1488 2912
rect 1552 2848 1748 2912
rect 1812 2848 2008 2912
rect 2072 2848 2268 2912
rect 2332 2848 2528 2912
rect 2592 2848 2788 2912
rect 2852 2848 3048 2912
rect 3112 2848 3308 2912
rect 3372 2848 3568 2912
rect 3632 2848 3828 2912
rect 3892 2848 4088 2912
rect 4152 2848 4348 2912
rect 4412 2848 4608 2912
rect 4672 2848 4868 2912
rect 4932 2848 5128 2912
rect 5192 2848 5470 2912
rect -770 2830 5470 2848
rect 6030 -2460 6130 -2360
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_0
timestamp 1757161594
transform 0 1 3007 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_1
timestamp 1757161594
transform 0 1 2227 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_2
timestamp 1757161594
transform 0 1 407 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_3
timestamp 1757161594
transform 0 1 2487 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_4
timestamp 1757161594
transform 0 1 927 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_5
timestamp 1757161594
transform 0 1 667 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_6
timestamp 1757161594
transform 0 1 147 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_7
timestamp 1757161594
transform 0 1 2747 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_8
timestamp 1757161594
transform 0 1 1447 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_9
timestamp 1757161594
transform 0 1 1187 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_10
timestamp 1757161594
transform 0 1 1707 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_11
timestamp 1757161594
transform 0 1 1967 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_12
timestamp 1757161594
transform 0 1 5347 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_13
timestamp 1757161594
transform 0 1 -113 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_14
timestamp 1757161594
transform 0 1 147 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_16
timestamp 1757161594
transform 0 1 3267 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_17
timestamp 1757161594
transform 0 1 3527 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_18
timestamp 1757161594
transform 0 1 3787 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_19
timestamp 1757161594
transform 0 1 4047 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_20
timestamp 1757161594
transform 0 1 4307 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_21
timestamp 1757161594
transform 0 1 4567 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_22
timestamp 1757161594
transform 0 1 4827 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_23
timestamp 1757161594
transform 0 1 5087 -1 0 1148
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_24
timestamp 1757161594
transform 0 1 1447 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_25
timestamp 1757161594
transform 0 1 1707 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_26
timestamp 1757161594
transform 0 1 927 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_27
timestamp 1757161594
transform 0 1 1187 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_28
timestamp 1757161594
transform 0 1 407 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_29
timestamp 1757161594
transform 0 1 667 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_30
timestamp 1757161594
transform 0 1 3007 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_31
timestamp 1757161594
transform 0 1 3267 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_32
timestamp 1757161594
transform 0 1 3527 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_33
timestamp 1757161594
transform 0 1 2747 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_34
timestamp 1757161594
transform 0 1 1967 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_35
timestamp 1757161594
transform 0 1 2227 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_36
timestamp 1757161594
transform 0 1 2487 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_37
timestamp 1757161594
transform 0 1 4827 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_38
timestamp 1757161594
transform 0 1 5087 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_39
timestamp 1757161594
transform 0 1 4307 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_40
timestamp 1757161594
transform 0 1 4567 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_41
timestamp 1757161594
transform 0 1 3787 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_42
timestamp 1757161594
transform 0 1 4047 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_43
timestamp 1757161594
transform 0 1 5347 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_G235U9  sky130_fd_pr__nfet_01v8_lvt_G235U9_44
timestamp 1757161594
transform 0 1 -113 -1 0 -1182
box -1084 -107 1084 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_0
timestamp 1757161594
transform 0 1 147 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_1
timestamp 1757161594
transform 0 1 -113 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_2
timestamp 1757161594
transform 0 1 1707 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_3
timestamp 1757161594
transform 0 1 407 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_4
timestamp 1757161594
transform 0 1 667 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_5
timestamp 1757161594
transform 0 1 927 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_6
timestamp 1757161594
transform 0 1 1447 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_7
timestamp 1757161594
transform 0 1 1187 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_9
timestamp 1757161594
transform 0 1 2487 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_10
timestamp 1757161594
transform 0 1 2747 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_11
timestamp 1757161594
transform 0 1 3007 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_12
timestamp 1757161594
transform 0 1 3267 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_13
timestamp 1757161594
transform 0 1 3527 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_14
timestamp 1757161594
transform 0 1 1967 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_15
timestamp 1757161594
transform 0 1 3787 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_16
timestamp 1757161594
transform 0 1 4047 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_17
timestamp 1757161594
transform 0 1 4307 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_18
timestamp 1757161594
transform 0 1 4567 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_19
timestamp 1757161594
transform 0 1 4827 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_20
timestamp 1757161594
transform 0 1 5087 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_21
timestamp 1757161594
transform 0 1 5347 -1 0 -2562
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_22
timestamp 1757161594
transform 0 1 667 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_23
timestamp 1757161594
transform 0 1 407 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_24
timestamp 1757161594
transform 0 1 147 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_25
timestamp 1757161594
transform 0 1 -113 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_26
timestamp 1757161594
transform 0 1 2487 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_27
timestamp 1757161594
transform 0 1 2747 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_28
timestamp 1757161594
transform 0 1 3007 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_29
timestamp 1757161594
transform 0 1 1707 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_30
timestamp 1757161594
transform 0 1 1967 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_31
timestamp 1757161594
transform 0 1 2227 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_32
timestamp 1757161594
transform 0 1 927 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_33
timestamp 1757161594
transform 0 1 1187 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_34
timestamp 1757161594
transform 0 1 1447 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_35
timestamp 1757161594
transform 0 1 4827 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_36
timestamp 1757161594
transform 0 1 5087 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_37
timestamp 1757161594
transform 0 1 5347 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_38
timestamp 1757161594
transform 0 1 4047 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_39
timestamp 1757161594
transform 0 1 4307 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_40
timestamp 1757161594
transform 0 1 4567 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_41
timestamp 1757161594
transform 0 1 3267 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_42
timestamp 1757161594
transform 0 1 3527 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_43
timestamp 1757161594
transform 0 1 3787 -1 0 2518
box -134 -107 134 107
use sky130_fd_pr__nfet_01v8_lvt_QGGREF  sky130_fd_pr__nfet_01v8_lvt_QGGREF_44
timestamp 1757161594
transform 0 1 2227 -1 0 -2562
box -134 -107 134 107
<< labels >>
flabel metal4 s -770 2830 -680 2930 0 FreeSans 782 0 0 0 Vbias1
port 0 nsew
<< end >>
