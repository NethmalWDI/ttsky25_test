magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -163 8977 6143 9063
rect -163 -107 -77 8977
rect 6057 -107 6143 8977
rect -163 -193 6143 -107
<< psubdiff >>
rect -137 9003 -33 9037
rect 1 9003 35 9037
rect 69 9003 103 9037
rect 137 9003 171 9037
rect 205 9003 239 9037
rect 273 9003 307 9037
rect 341 9003 375 9037
rect 409 9003 443 9037
rect 477 9003 511 9037
rect 545 9003 579 9037
rect 613 9003 647 9037
rect 681 9003 715 9037
rect 749 9003 783 9037
rect 817 9003 851 9037
rect 885 9003 919 9037
rect 953 9003 987 9037
rect 1021 9003 1055 9037
rect 1089 9003 1123 9037
rect 1157 9003 1191 9037
rect 1225 9003 1259 9037
rect 1293 9003 1327 9037
rect 1361 9003 1395 9037
rect 1429 9003 1463 9037
rect 1497 9003 1531 9037
rect 1565 9003 1599 9037
rect 1633 9003 1667 9037
rect 1701 9003 1735 9037
rect 1769 9003 1803 9037
rect 1837 9003 1871 9037
rect 1905 9003 1939 9037
rect 1973 9003 2007 9037
rect 2041 9003 2075 9037
rect 2109 9003 2143 9037
rect 2177 9003 2211 9037
rect 2245 9003 2279 9037
rect 2313 9003 2347 9037
rect 2381 9003 2415 9037
rect 2449 9003 2483 9037
rect 2517 9003 2551 9037
rect 2585 9003 2619 9037
rect 2653 9003 2687 9037
rect 2721 9003 2755 9037
rect 2789 9003 2823 9037
rect 2857 9003 2891 9037
rect 2925 9003 2959 9037
rect 2993 9003 3027 9037
rect 3061 9003 3095 9037
rect 3129 9003 3163 9037
rect 3197 9003 3231 9037
rect 3265 9003 3299 9037
rect 3333 9003 3367 9037
rect 3401 9003 3435 9037
rect 3469 9003 3503 9037
rect 3537 9003 3571 9037
rect 3605 9003 3639 9037
rect 3673 9003 3707 9037
rect 3741 9003 3775 9037
rect 3809 9003 3843 9037
rect 3877 9003 3911 9037
rect 3945 9003 3979 9037
rect 4013 9003 4047 9037
rect 4081 9003 4115 9037
rect 4149 9003 4183 9037
rect 4217 9003 4251 9037
rect 4285 9003 4319 9037
rect 4353 9003 4387 9037
rect 4421 9003 4455 9037
rect 4489 9003 4523 9037
rect 4557 9003 4591 9037
rect 4625 9003 4659 9037
rect 4693 9003 4727 9037
rect 4761 9003 4795 9037
rect 4829 9003 4863 9037
rect 4897 9003 4931 9037
rect 4965 9003 4999 9037
rect 5033 9003 5067 9037
rect 5101 9003 5135 9037
rect 5169 9003 5203 9037
rect 5237 9003 5271 9037
rect 5305 9003 5339 9037
rect 5373 9003 5407 9037
rect 5441 9003 5475 9037
rect 5509 9003 5543 9037
rect 5577 9003 5611 9037
rect 5645 9003 5679 9037
rect 5713 9003 5747 9037
rect 5781 9003 5815 9037
rect 5849 9003 5883 9037
rect 5917 9003 5951 9037
rect 5985 9003 6019 9037
rect 6053 9003 6117 9037
rect -137 8967 -103 9003
rect -137 8899 -103 8933
rect -137 8831 -103 8865
rect -137 8763 -103 8797
rect -137 8695 -103 8729
rect -137 8627 -103 8661
rect -137 8559 -103 8593
rect -137 8491 -103 8525
rect -137 8423 -103 8457
rect -137 8355 -103 8389
rect -137 8287 -103 8321
rect -137 8219 -103 8253
rect -137 8151 -103 8185
rect -137 8083 -103 8117
rect -137 8015 -103 8049
rect -137 7947 -103 7981
rect -137 7879 -103 7913
rect -137 7811 -103 7845
rect -137 7743 -103 7777
rect -137 7675 -103 7709
rect -137 7607 -103 7641
rect -137 7539 -103 7573
rect -137 7471 -103 7505
rect -137 7403 -103 7437
rect -137 7335 -103 7369
rect -137 7267 -103 7301
rect -137 7199 -103 7233
rect -137 7131 -103 7165
rect -137 7063 -103 7097
rect -137 6995 -103 7029
rect -137 6927 -103 6961
rect -137 6859 -103 6893
rect -137 6791 -103 6825
rect -137 6723 -103 6757
rect -137 6655 -103 6689
rect -137 6587 -103 6621
rect -137 6519 -103 6553
rect -137 6451 -103 6485
rect -137 6383 -103 6417
rect -137 6315 -103 6349
rect -137 6247 -103 6281
rect -137 6179 -103 6213
rect -137 6111 -103 6145
rect -137 6043 -103 6077
rect -137 5975 -103 6009
rect -137 5907 -103 5941
rect -137 5839 -103 5873
rect -137 5771 -103 5805
rect -137 5703 -103 5737
rect -137 5635 -103 5669
rect -137 5567 -103 5601
rect -137 5499 -103 5533
rect -137 5431 -103 5465
rect -137 5363 -103 5397
rect -137 5295 -103 5329
rect -137 5227 -103 5261
rect -137 5159 -103 5193
rect -137 5091 -103 5125
rect -137 5023 -103 5057
rect -137 4955 -103 4989
rect -137 4887 -103 4921
rect -137 4819 -103 4853
rect -137 4751 -103 4785
rect -137 4683 -103 4717
rect -137 4615 -103 4649
rect -137 4547 -103 4581
rect -137 4479 -103 4513
rect -137 4411 -103 4445
rect -137 4343 -103 4377
rect -137 4275 -103 4309
rect -137 4207 -103 4241
rect -137 4139 -103 4173
rect -137 4071 -103 4105
rect -137 4003 -103 4037
rect -137 3935 -103 3969
rect -137 3867 -103 3901
rect -137 3799 -103 3833
rect -137 3731 -103 3765
rect -137 3663 -103 3697
rect -137 3595 -103 3629
rect -137 3527 -103 3561
rect -137 3459 -103 3493
rect -137 3391 -103 3425
rect -137 3323 -103 3357
rect -137 3255 -103 3289
rect -137 3187 -103 3221
rect -137 3119 -103 3153
rect -137 3051 -103 3085
rect -137 2983 -103 3017
rect -137 2915 -103 2949
rect -137 2847 -103 2881
rect -137 2779 -103 2813
rect -137 2711 -103 2745
rect -137 2643 -103 2677
rect -137 2575 -103 2609
rect -137 2507 -103 2541
rect -137 2439 -103 2473
rect -137 2371 -103 2405
rect -137 2303 -103 2337
rect -137 2235 -103 2269
rect -137 2167 -103 2201
rect -137 2099 -103 2133
rect -137 2031 -103 2065
rect -137 1963 -103 1997
rect -137 1895 -103 1929
rect -137 1827 -103 1861
rect -137 1759 -103 1793
rect -137 1691 -103 1725
rect -137 1623 -103 1657
rect -137 1555 -103 1589
rect -137 1487 -103 1521
rect -137 1419 -103 1453
rect -137 1351 -103 1385
rect -137 1283 -103 1317
rect -137 1215 -103 1249
rect -137 1147 -103 1181
rect -137 1079 -103 1113
rect -137 1011 -103 1045
rect -137 943 -103 977
rect -137 875 -103 909
rect -137 807 -103 841
rect -137 739 -103 773
rect -137 671 -103 705
rect -137 603 -103 637
rect -137 535 -103 569
rect -137 467 -103 501
rect -137 399 -103 433
rect -137 331 -103 365
rect -137 263 -103 297
rect -137 195 -103 229
rect -137 127 -103 161
rect -137 59 -103 93
rect -137 -9 -103 25
rect -137 -77 -103 -43
rect -137 -133 -103 -111
rect 6083 8974 6117 9003
rect 6083 8906 6117 8940
rect 6083 8838 6117 8872
rect 6083 8770 6117 8804
rect 6083 8702 6117 8736
rect 6083 8634 6117 8668
rect 6083 8566 6117 8600
rect 6083 8498 6117 8532
rect 6083 8430 6117 8464
rect 6083 8362 6117 8396
rect 6083 8294 6117 8328
rect 6083 8226 6117 8260
rect 6083 8158 6117 8192
rect 6083 8090 6117 8124
rect 6083 8022 6117 8056
rect 6083 7954 6117 7988
rect 6083 7886 6117 7920
rect 6083 7818 6117 7852
rect 6083 7750 6117 7784
rect 6083 7682 6117 7716
rect 6083 7614 6117 7648
rect 6083 7546 6117 7580
rect 6083 7478 6117 7512
rect 6083 7410 6117 7444
rect 6083 7342 6117 7376
rect 6083 7274 6117 7308
rect 6083 7206 6117 7240
rect 6083 7138 6117 7172
rect 6083 7070 6117 7104
rect 6083 7002 6117 7036
rect 6083 6934 6117 6968
rect 6083 6866 6117 6900
rect 6083 6798 6117 6832
rect 6083 6730 6117 6764
rect 6083 6662 6117 6696
rect 6083 6594 6117 6628
rect 6083 6526 6117 6560
rect 6083 6458 6117 6492
rect 6083 6390 6117 6424
rect 6083 6322 6117 6356
rect 6083 6254 6117 6288
rect 6083 6186 6117 6220
rect 6083 6118 6117 6152
rect 6083 6050 6117 6084
rect 6083 5982 6117 6016
rect 6083 5914 6117 5948
rect 6083 5846 6117 5880
rect 6083 5778 6117 5812
rect 6083 5710 6117 5744
rect 6083 5642 6117 5676
rect 6083 5574 6117 5608
rect 6083 5506 6117 5540
rect 6083 5438 6117 5472
rect 6083 5370 6117 5404
rect 6083 5302 6117 5336
rect 6083 5234 6117 5268
rect 6083 5166 6117 5200
rect 6083 5098 6117 5132
rect 6083 5030 6117 5064
rect 6083 4962 6117 4996
rect 6083 4894 6117 4928
rect 6083 4826 6117 4860
rect 6083 4758 6117 4792
rect 6083 4690 6117 4724
rect 6083 4622 6117 4656
rect 6083 4554 6117 4588
rect 6083 4486 6117 4520
rect 6083 4418 6117 4452
rect 6083 4350 6117 4384
rect 6083 4282 6117 4316
rect 6083 4214 6117 4248
rect 6083 4146 6117 4180
rect 6083 4078 6117 4112
rect 6083 4010 6117 4044
rect 6083 3942 6117 3976
rect 6083 3874 6117 3908
rect 6083 3806 6117 3840
rect 6083 3738 6117 3772
rect 6083 3670 6117 3704
rect 6083 3602 6117 3636
rect 6083 3534 6117 3568
rect 6083 3466 6117 3500
rect 6083 3398 6117 3432
rect 6083 3330 6117 3364
rect 6083 3262 6117 3296
rect 6083 3194 6117 3228
rect 6083 3126 6117 3160
rect 6083 3058 6117 3092
rect 6083 2990 6117 3024
rect 6083 2922 6117 2956
rect 6083 2854 6117 2888
rect 6083 2786 6117 2820
rect 6083 2718 6117 2752
rect 6083 2650 6117 2684
rect 6083 2582 6117 2616
rect 6083 2514 6117 2548
rect 6083 2446 6117 2480
rect 6083 2378 6117 2412
rect 6083 2310 6117 2344
rect 6083 2242 6117 2276
rect 6083 2174 6117 2208
rect 6083 2106 6117 2140
rect 6083 2038 6117 2072
rect 6083 1970 6117 2004
rect 6083 1902 6117 1936
rect 6083 1834 6117 1868
rect 6083 1766 6117 1800
rect 6083 1698 6117 1732
rect 6083 1630 6117 1664
rect 6083 1562 6117 1596
rect 6083 1494 6117 1528
rect 6083 1426 6117 1460
rect 6083 1358 6117 1392
rect 6083 1290 6117 1324
rect 6083 1222 6117 1256
rect 6083 1154 6117 1188
rect 6083 1086 6117 1120
rect 6083 1018 6117 1052
rect 6083 950 6117 984
rect 6083 882 6117 916
rect 6083 814 6117 848
rect 6083 746 6117 780
rect 6083 678 6117 712
rect 6083 610 6117 644
rect 6083 542 6117 576
rect 6083 474 6117 508
rect 6083 406 6117 440
rect 6083 338 6117 372
rect 6083 270 6117 304
rect 6083 202 6117 236
rect 6083 134 6117 168
rect 6083 66 6117 100
rect 6083 -2 6117 32
rect 6083 -70 6117 -36
rect 6083 -133 6117 -104
rect -137 -167 -33 -133
rect 1 -167 35 -133
rect 69 -167 103 -133
rect 137 -167 171 -133
rect 205 -167 239 -133
rect 273 -167 307 -133
rect 341 -167 375 -133
rect 409 -167 443 -133
rect 477 -167 511 -133
rect 545 -167 579 -133
rect 613 -167 647 -133
rect 681 -167 715 -133
rect 749 -167 783 -133
rect 817 -167 851 -133
rect 885 -167 919 -133
rect 953 -167 987 -133
rect 1021 -167 1055 -133
rect 1089 -167 1123 -133
rect 1157 -167 1191 -133
rect 1225 -167 1259 -133
rect 1293 -167 1327 -133
rect 1361 -167 1395 -133
rect 1429 -167 1463 -133
rect 1497 -167 1531 -133
rect 1565 -167 1599 -133
rect 1633 -167 1667 -133
rect 1701 -167 1735 -133
rect 1769 -167 1803 -133
rect 1837 -167 1871 -133
rect 1905 -167 1939 -133
rect 1973 -167 2007 -133
rect 2041 -167 2075 -133
rect 2109 -167 2143 -133
rect 2177 -167 2211 -133
rect 2245 -167 2279 -133
rect 2313 -167 2347 -133
rect 2381 -167 2415 -133
rect 2449 -167 2483 -133
rect 2517 -167 2551 -133
rect 2585 -167 2619 -133
rect 2653 -167 2687 -133
rect 2721 -167 2755 -133
rect 2789 -167 2823 -133
rect 2857 -167 2891 -133
rect 2925 -167 2959 -133
rect 2993 -167 3027 -133
rect 3061 -167 3095 -133
rect 3129 -167 3163 -133
rect 3197 -167 3231 -133
rect 3265 -167 3299 -133
rect 3333 -167 3367 -133
rect 3401 -167 3435 -133
rect 3469 -167 3503 -133
rect 3537 -167 3571 -133
rect 3605 -167 3639 -133
rect 3673 -167 3707 -133
rect 3741 -167 3775 -133
rect 3809 -167 3843 -133
rect 3877 -167 3911 -133
rect 3945 -167 3979 -133
rect 4013 -167 4047 -133
rect 4081 -167 4115 -133
rect 4149 -167 4183 -133
rect 4217 -167 4251 -133
rect 4285 -167 4319 -133
rect 4353 -167 4387 -133
rect 4421 -167 4455 -133
rect 4489 -167 4523 -133
rect 4557 -167 4591 -133
rect 4625 -167 4659 -133
rect 4693 -167 4727 -133
rect 4761 -167 4795 -133
rect 4829 -167 4863 -133
rect 4897 -167 4931 -133
rect 4965 -167 4999 -133
rect 5033 -167 5067 -133
rect 5101 -167 5135 -133
rect 5169 -167 5203 -133
rect 5237 -167 5271 -133
rect 5305 -167 5339 -133
rect 5373 -167 5407 -133
rect 5441 -167 5475 -133
rect 5509 -167 5543 -133
rect 5577 -167 5611 -133
rect 5645 -167 5679 -133
rect 5713 -167 5747 -133
rect 5781 -167 5815 -133
rect 5849 -167 5883 -133
rect 5917 -167 5951 -133
rect 5985 -167 6019 -133
rect 6053 -167 6117 -133
<< psubdiffcont >>
rect -33 9003 1 9037
rect 35 9003 69 9037
rect 103 9003 137 9037
rect 171 9003 205 9037
rect 239 9003 273 9037
rect 307 9003 341 9037
rect 375 9003 409 9037
rect 443 9003 477 9037
rect 511 9003 545 9037
rect 579 9003 613 9037
rect 647 9003 681 9037
rect 715 9003 749 9037
rect 783 9003 817 9037
rect 851 9003 885 9037
rect 919 9003 953 9037
rect 987 9003 1021 9037
rect 1055 9003 1089 9037
rect 1123 9003 1157 9037
rect 1191 9003 1225 9037
rect 1259 9003 1293 9037
rect 1327 9003 1361 9037
rect 1395 9003 1429 9037
rect 1463 9003 1497 9037
rect 1531 9003 1565 9037
rect 1599 9003 1633 9037
rect 1667 9003 1701 9037
rect 1735 9003 1769 9037
rect 1803 9003 1837 9037
rect 1871 9003 1905 9037
rect 1939 9003 1973 9037
rect 2007 9003 2041 9037
rect 2075 9003 2109 9037
rect 2143 9003 2177 9037
rect 2211 9003 2245 9037
rect 2279 9003 2313 9037
rect 2347 9003 2381 9037
rect 2415 9003 2449 9037
rect 2483 9003 2517 9037
rect 2551 9003 2585 9037
rect 2619 9003 2653 9037
rect 2687 9003 2721 9037
rect 2755 9003 2789 9037
rect 2823 9003 2857 9037
rect 2891 9003 2925 9037
rect 2959 9003 2993 9037
rect 3027 9003 3061 9037
rect 3095 9003 3129 9037
rect 3163 9003 3197 9037
rect 3231 9003 3265 9037
rect 3299 9003 3333 9037
rect 3367 9003 3401 9037
rect 3435 9003 3469 9037
rect 3503 9003 3537 9037
rect 3571 9003 3605 9037
rect 3639 9003 3673 9037
rect 3707 9003 3741 9037
rect 3775 9003 3809 9037
rect 3843 9003 3877 9037
rect 3911 9003 3945 9037
rect 3979 9003 4013 9037
rect 4047 9003 4081 9037
rect 4115 9003 4149 9037
rect 4183 9003 4217 9037
rect 4251 9003 4285 9037
rect 4319 9003 4353 9037
rect 4387 9003 4421 9037
rect 4455 9003 4489 9037
rect 4523 9003 4557 9037
rect 4591 9003 4625 9037
rect 4659 9003 4693 9037
rect 4727 9003 4761 9037
rect 4795 9003 4829 9037
rect 4863 9003 4897 9037
rect 4931 9003 4965 9037
rect 4999 9003 5033 9037
rect 5067 9003 5101 9037
rect 5135 9003 5169 9037
rect 5203 9003 5237 9037
rect 5271 9003 5305 9037
rect 5339 9003 5373 9037
rect 5407 9003 5441 9037
rect 5475 9003 5509 9037
rect 5543 9003 5577 9037
rect 5611 9003 5645 9037
rect 5679 9003 5713 9037
rect 5747 9003 5781 9037
rect 5815 9003 5849 9037
rect 5883 9003 5917 9037
rect 5951 9003 5985 9037
rect 6019 9003 6053 9037
rect -137 8933 -103 8967
rect -137 8865 -103 8899
rect -137 8797 -103 8831
rect -137 8729 -103 8763
rect -137 8661 -103 8695
rect -137 8593 -103 8627
rect -137 8525 -103 8559
rect -137 8457 -103 8491
rect -137 8389 -103 8423
rect -137 8321 -103 8355
rect -137 8253 -103 8287
rect -137 8185 -103 8219
rect -137 8117 -103 8151
rect -137 8049 -103 8083
rect -137 7981 -103 8015
rect -137 7913 -103 7947
rect -137 7845 -103 7879
rect -137 7777 -103 7811
rect -137 7709 -103 7743
rect -137 7641 -103 7675
rect -137 7573 -103 7607
rect -137 7505 -103 7539
rect -137 7437 -103 7471
rect -137 7369 -103 7403
rect -137 7301 -103 7335
rect -137 7233 -103 7267
rect -137 7165 -103 7199
rect -137 7097 -103 7131
rect -137 7029 -103 7063
rect -137 6961 -103 6995
rect -137 6893 -103 6927
rect -137 6825 -103 6859
rect -137 6757 -103 6791
rect -137 6689 -103 6723
rect -137 6621 -103 6655
rect -137 6553 -103 6587
rect -137 6485 -103 6519
rect -137 6417 -103 6451
rect -137 6349 -103 6383
rect -137 6281 -103 6315
rect -137 6213 -103 6247
rect -137 6145 -103 6179
rect -137 6077 -103 6111
rect -137 6009 -103 6043
rect -137 5941 -103 5975
rect -137 5873 -103 5907
rect -137 5805 -103 5839
rect -137 5737 -103 5771
rect -137 5669 -103 5703
rect -137 5601 -103 5635
rect -137 5533 -103 5567
rect -137 5465 -103 5499
rect -137 5397 -103 5431
rect -137 5329 -103 5363
rect -137 5261 -103 5295
rect -137 5193 -103 5227
rect -137 5125 -103 5159
rect -137 5057 -103 5091
rect -137 4989 -103 5023
rect -137 4921 -103 4955
rect -137 4853 -103 4887
rect -137 4785 -103 4819
rect -137 4717 -103 4751
rect -137 4649 -103 4683
rect -137 4581 -103 4615
rect -137 4513 -103 4547
rect -137 4445 -103 4479
rect -137 4377 -103 4411
rect -137 4309 -103 4343
rect -137 4241 -103 4275
rect -137 4173 -103 4207
rect -137 4105 -103 4139
rect -137 4037 -103 4071
rect -137 3969 -103 4003
rect -137 3901 -103 3935
rect -137 3833 -103 3867
rect -137 3765 -103 3799
rect -137 3697 -103 3731
rect -137 3629 -103 3663
rect -137 3561 -103 3595
rect -137 3493 -103 3527
rect -137 3425 -103 3459
rect -137 3357 -103 3391
rect -137 3289 -103 3323
rect -137 3221 -103 3255
rect -137 3153 -103 3187
rect -137 3085 -103 3119
rect -137 3017 -103 3051
rect -137 2949 -103 2983
rect -137 2881 -103 2915
rect -137 2813 -103 2847
rect -137 2745 -103 2779
rect -137 2677 -103 2711
rect -137 2609 -103 2643
rect -137 2541 -103 2575
rect -137 2473 -103 2507
rect -137 2405 -103 2439
rect -137 2337 -103 2371
rect -137 2269 -103 2303
rect -137 2201 -103 2235
rect -137 2133 -103 2167
rect -137 2065 -103 2099
rect -137 1997 -103 2031
rect -137 1929 -103 1963
rect -137 1861 -103 1895
rect -137 1793 -103 1827
rect -137 1725 -103 1759
rect -137 1657 -103 1691
rect -137 1589 -103 1623
rect -137 1521 -103 1555
rect -137 1453 -103 1487
rect -137 1385 -103 1419
rect -137 1317 -103 1351
rect -137 1249 -103 1283
rect -137 1181 -103 1215
rect -137 1113 -103 1147
rect -137 1045 -103 1079
rect -137 977 -103 1011
rect -137 909 -103 943
rect -137 841 -103 875
rect -137 773 -103 807
rect -137 705 -103 739
rect -137 637 -103 671
rect -137 569 -103 603
rect -137 501 -103 535
rect -137 433 -103 467
rect -137 365 -103 399
rect -137 297 -103 331
rect -137 229 -103 263
rect -137 161 -103 195
rect -137 93 -103 127
rect -137 25 -103 59
rect -137 -43 -103 -9
rect -137 -111 -103 -77
rect 6083 8940 6117 8974
rect 6083 8872 6117 8906
rect 6083 8804 6117 8838
rect 6083 8736 6117 8770
rect 6083 8668 6117 8702
rect 6083 8600 6117 8634
rect 6083 8532 6117 8566
rect 6083 8464 6117 8498
rect 6083 8396 6117 8430
rect 6083 8328 6117 8362
rect 6083 8260 6117 8294
rect 6083 8192 6117 8226
rect 6083 8124 6117 8158
rect 6083 8056 6117 8090
rect 6083 7988 6117 8022
rect 6083 7920 6117 7954
rect 6083 7852 6117 7886
rect 6083 7784 6117 7818
rect 6083 7716 6117 7750
rect 6083 7648 6117 7682
rect 6083 7580 6117 7614
rect 6083 7512 6117 7546
rect 6083 7444 6117 7478
rect 6083 7376 6117 7410
rect 6083 7308 6117 7342
rect 6083 7240 6117 7274
rect 6083 7172 6117 7206
rect 6083 7104 6117 7138
rect 6083 7036 6117 7070
rect 6083 6968 6117 7002
rect 6083 6900 6117 6934
rect 6083 6832 6117 6866
rect 6083 6764 6117 6798
rect 6083 6696 6117 6730
rect 6083 6628 6117 6662
rect 6083 6560 6117 6594
rect 6083 6492 6117 6526
rect 6083 6424 6117 6458
rect 6083 6356 6117 6390
rect 6083 6288 6117 6322
rect 6083 6220 6117 6254
rect 6083 6152 6117 6186
rect 6083 6084 6117 6118
rect 6083 6016 6117 6050
rect 6083 5948 6117 5982
rect 6083 5880 6117 5914
rect 6083 5812 6117 5846
rect 6083 5744 6117 5778
rect 6083 5676 6117 5710
rect 6083 5608 6117 5642
rect 6083 5540 6117 5574
rect 6083 5472 6117 5506
rect 6083 5404 6117 5438
rect 6083 5336 6117 5370
rect 6083 5268 6117 5302
rect 6083 5200 6117 5234
rect 6083 5132 6117 5166
rect 6083 5064 6117 5098
rect 6083 4996 6117 5030
rect 6083 4928 6117 4962
rect 6083 4860 6117 4894
rect 6083 4792 6117 4826
rect 6083 4724 6117 4758
rect 6083 4656 6117 4690
rect 6083 4588 6117 4622
rect 6083 4520 6117 4554
rect 6083 4452 6117 4486
rect 6083 4384 6117 4418
rect 6083 4316 6117 4350
rect 6083 4248 6117 4282
rect 6083 4180 6117 4214
rect 6083 4112 6117 4146
rect 6083 4044 6117 4078
rect 6083 3976 6117 4010
rect 6083 3908 6117 3942
rect 6083 3840 6117 3874
rect 6083 3772 6117 3806
rect 6083 3704 6117 3738
rect 6083 3636 6117 3670
rect 6083 3568 6117 3602
rect 6083 3500 6117 3534
rect 6083 3432 6117 3466
rect 6083 3364 6117 3398
rect 6083 3296 6117 3330
rect 6083 3228 6117 3262
rect 6083 3160 6117 3194
rect 6083 3092 6117 3126
rect 6083 3024 6117 3058
rect 6083 2956 6117 2990
rect 6083 2888 6117 2922
rect 6083 2820 6117 2854
rect 6083 2752 6117 2786
rect 6083 2684 6117 2718
rect 6083 2616 6117 2650
rect 6083 2548 6117 2582
rect 6083 2480 6117 2514
rect 6083 2412 6117 2446
rect 6083 2344 6117 2378
rect 6083 2276 6117 2310
rect 6083 2208 6117 2242
rect 6083 2140 6117 2174
rect 6083 2072 6117 2106
rect 6083 2004 6117 2038
rect 6083 1936 6117 1970
rect 6083 1868 6117 1902
rect 6083 1800 6117 1834
rect 6083 1732 6117 1766
rect 6083 1664 6117 1698
rect 6083 1596 6117 1630
rect 6083 1528 6117 1562
rect 6083 1460 6117 1494
rect 6083 1392 6117 1426
rect 6083 1324 6117 1358
rect 6083 1256 6117 1290
rect 6083 1188 6117 1222
rect 6083 1120 6117 1154
rect 6083 1052 6117 1086
rect 6083 984 6117 1018
rect 6083 916 6117 950
rect 6083 848 6117 882
rect 6083 780 6117 814
rect 6083 712 6117 746
rect 6083 644 6117 678
rect 6083 576 6117 610
rect 6083 508 6117 542
rect 6083 440 6117 474
rect 6083 372 6117 406
rect 6083 304 6117 338
rect 6083 236 6117 270
rect 6083 168 6117 202
rect 6083 100 6117 134
rect 6083 32 6117 66
rect 6083 -36 6117 -2
rect 6083 -104 6117 -70
rect -33 -167 1 -133
rect 35 -167 69 -133
rect 103 -167 137 -133
rect 171 -167 205 -133
rect 239 -167 273 -133
rect 307 -167 341 -133
rect 375 -167 409 -133
rect 443 -167 477 -133
rect 511 -167 545 -133
rect 579 -167 613 -133
rect 647 -167 681 -133
rect 715 -167 749 -133
rect 783 -167 817 -133
rect 851 -167 885 -133
rect 919 -167 953 -133
rect 987 -167 1021 -133
rect 1055 -167 1089 -133
rect 1123 -167 1157 -133
rect 1191 -167 1225 -133
rect 1259 -167 1293 -133
rect 1327 -167 1361 -133
rect 1395 -167 1429 -133
rect 1463 -167 1497 -133
rect 1531 -167 1565 -133
rect 1599 -167 1633 -133
rect 1667 -167 1701 -133
rect 1735 -167 1769 -133
rect 1803 -167 1837 -133
rect 1871 -167 1905 -133
rect 1939 -167 1973 -133
rect 2007 -167 2041 -133
rect 2075 -167 2109 -133
rect 2143 -167 2177 -133
rect 2211 -167 2245 -133
rect 2279 -167 2313 -133
rect 2347 -167 2381 -133
rect 2415 -167 2449 -133
rect 2483 -167 2517 -133
rect 2551 -167 2585 -133
rect 2619 -167 2653 -133
rect 2687 -167 2721 -133
rect 2755 -167 2789 -133
rect 2823 -167 2857 -133
rect 2891 -167 2925 -133
rect 2959 -167 2993 -133
rect 3027 -167 3061 -133
rect 3095 -167 3129 -133
rect 3163 -167 3197 -133
rect 3231 -167 3265 -133
rect 3299 -167 3333 -133
rect 3367 -167 3401 -133
rect 3435 -167 3469 -133
rect 3503 -167 3537 -133
rect 3571 -167 3605 -133
rect 3639 -167 3673 -133
rect 3707 -167 3741 -133
rect 3775 -167 3809 -133
rect 3843 -167 3877 -133
rect 3911 -167 3945 -133
rect 3979 -167 4013 -133
rect 4047 -167 4081 -133
rect 4115 -167 4149 -133
rect 4183 -167 4217 -133
rect 4251 -167 4285 -133
rect 4319 -167 4353 -133
rect 4387 -167 4421 -133
rect 4455 -167 4489 -133
rect 4523 -167 4557 -133
rect 4591 -167 4625 -133
rect 4659 -167 4693 -133
rect 4727 -167 4761 -133
rect 4795 -167 4829 -133
rect 4863 -167 4897 -133
rect 4931 -167 4965 -133
rect 4999 -167 5033 -133
rect 5067 -167 5101 -133
rect 5135 -167 5169 -133
rect 5203 -167 5237 -133
rect 5271 -167 5305 -133
rect 5339 -167 5373 -133
rect 5407 -167 5441 -133
rect 5475 -167 5509 -133
rect 5543 -167 5577 -133
rect 5611 -167 5645 -133
rect 5679 -167 5713 -133
rect 5747 -167 5781 -133
rect 5815 -167 5849 -133
rect 5883 -167 5917 -133
rect 5951 -167 5985 -133
rect 6019 -167 6053 -133
<< locali >>
rect -137 9003 -33 9037
rect 1 9003 35 9037
rect 69 9003 103 9037
rect 137 9003 171 9037
rect 205 9003 239 9037
rect 273 9003 307 9037
rect 341 9003 375 9037
rect 409 9003 443 9037
rect 477 9003 511 9037
rect 545 9003 579 9037
rect 613 9003 647 9037
rect 681 9003 715 9037
rect 749 9003 783 9037
rect 817 9003 851 9037
rect 885 9003 919 9037
rect 953 9003 987 9037
rect 1021 9003 1055 9037
rect 1089 9003 1123 9037
rect 1157 9003 1191 9037
rect 1225 9003 1259 9037
rect 1293 9003 1327 9037
rect 1361 9003 1395 9037
rect 1429 9003 1463 9037
rect 1497 9003 1531 9037
rect 1565 9003 1599 9037
rect 1633 9003 1667 9037
rect 1701 9003 1735 9037
rect 1769 9003 1803 9037
rect 1837 9003 1871 9037
rect 1905 9003 1939 9037
rect 1973 9003 2007 9037
rect 2041 9003 2075 9037
rect 2109 9003 2143 9037
rect 2177 9003 2211 9037
rect 2245 9003 2279 9037
rect 2313 9003 2347 9037
rect 2381 9003 2415 9037
rect 2449 9003 2483 9037
rect 2517 9003 2551 9037
rect 2585 9003 2619 9037
rect 2653 9003 2687 9037
rect 2721 9003 2755 9037
rect 2789 9003 2823 9037
rect 2857 9003 2891 9037
rect 2925 9003 2959 9037
rect 2993 9003 3027 9037
rect 3061 9003 3095 9037
rect 3129 9003 3163 9037
rect 3197 9003 3231 9037
rect 3265 9003 3299 9037
rect 3333 9003 3367 9037
rect 3401 9003 3435 9037
rect 3469 9003 3503 9037
rect 3537 9003 3571 9037
rect 3605 9003 3639 9037
rect 3673 9003 3707 9037
rect 3741 9003 3775 9037
rect 3809 9003 3843 9037
rect 3877 9003 3911 9037
rect 3945 9003 3979 9037
rect 4013 9003 4047 9037
rect 4081 9003 4115 9037
rect 4149 9003 4183 9037
rect 4217 9003 4251 9037
rect 4285 9003 4319 9037
rect 4353 9003 4387 9037
rect 4421 9003 4455 9037
rect 4489 9003 4523 9037
rect 4557 9003 4591 9037
rect 4625 9003 4659 9037
rect 4693 9003 4727 9037
rect 4761 9003 4795 9037
rect 4829 9003 4863 9037
rect 4897 9003 4931 9037
rect 4965 9003 4999 9037
rect 5033 9003 5067 9037
rect 5101 9003 5135 9037
rect 5169 9003 5203 9037
rect 5237 9003 5271 9037
rect 5305 9003 5339 9037
rect 5373 9003 5407 9037
rect 5441 9003 5475 9037
rect 5509 9003 5543 9037
rect 5577 9003 5611 9037
rect 5645 9003 5679 9037
rect 5713 9003 5747 9037
rect 5781 9003 5815 9037
rect 5849 9003 5883 9037
rect 5917 9003 5951 9037
rect 5985 9003 6019 9037
rect 6053 9003 6117 9037
rect -137 8967 -103 9003
rect -137 8899 -103 8933
rect -137 8831 -103 8865
rect -137 8763 -103 8797
rect -137 8695 -103 8729
rect -137 8627 -103 8661
rect -137 8559 -103 8593
rect -137 8491 -103 8525
rect -137 8423 -103 8457
rect -137 8355 -103 8389
rect -137 8287 -103 8321
rect -137 8219 -103 8253
rect -137 8151 -103 8185
rect -137 8083 -103 8117
rect -137 8015 -103 8049
rect -137 7947 -103 7981
rect -137 7879 -103 7913
rect -137 7811 -103 7845
rect -137 7743 -103 7777
rect -137 7675 -103 7709
rect -137 7607 -103 7641
rect -137 7539 -103 7573
rect -137 7471 -103 7505
rect -137 7403 -103 7437
rect -137 7335 -103 7369
rect -137 7267 -103 7301
rect -137 7199 -103 7233
rect -137 7131 -103 7165
rect -137 7063 -103 7097
rect -137 6995 -103 7029
rect -137 6927 -103 6961
rect -137 6859 -103 6893
rect -137 6791 -103 6825
rect -137 6723 -103 6757
rect -137 6655 -103 6689
rect -137 6587 -103 6621
rect -137 6519 -103 6553
rect -137 6451 -103 6485
rect -137 6383 -103 6417
rect -137 6315 -103 6349
rect -137 6247 -103 6281
rect -137 6179 -103 6213
rect -137 6111 -103 6145
rect -137 6043 -103 6077
rect -137 5975 -103 6009
rect -137 5907 -103 5941
rect -137 5839 -103 5873
rect -137 5771 -103 5805
rect -137 5703 -103 5737
rect -137 5635 -103 5669
rect -137 5567 -103 5601
rect -137 5499 -103 5533
rect -137 5431 -103 5465
rect -137 5363 -103 5397
rect -137 5295 -103 5329
rect -137 5227 -103 5261
rect -137 5159 -103 5193
rect -137 5091 -103 5125
rect -137 5023 -103 5057
rect -137 4955 -103 4989
rect -137 4887 -103 4921
rect -137 4819 -103 4853
rect -137 4751 -103 4785
rect -137 4683 -103 4717
rect -137 4615 -103 4649
rect -137 4547 -103 4581
rect -137 4479 -103 4513
rect -137 4411 -103 4445
rect -137 4343 -103 4377
rect -137 4275 -103 4309
rect -137 4207 -103 4241
rect -137 4139 -103 4173
rect -137 4071 -103 4105
rect -137 4003 -103 4037
rect -137 3935 -103 3969
rect -137 3867 -103 3901
rect -137 3799 -103 3833
rect -137 3731 -103 3765
rect -137 3663 -103 3697
rect -137 3595 -103 3629
rect -137 3527 -103 3561
rect -137 3459 -103 3493
rect -137 3391 -103 3425
rect -137 3323 -103 3357
rect -137 3255 -103 3289
rect -137 3187 -103 3221
rect -137 3119 -103 3153
rect -137 3051 -103 3085
rect -137 2983 -103 3017
rect -137 2915 -103 2949
rect -137 2847 -103 2881
rect -137 2779 -103 2813
rect -137 2711 -103 2745
rect -137 2643 -103 2677
rect -137 2575 -103 2609
rect -137 2507 -103 2541
rect -137 2439 -103 2473
rect -137 2371 -103 2405
rect -137 2303 -103 2337
rect -137 2235 -103 2269
rect -137 2167 -103 2201
rect -137 2099 -103 2133
rect -137 2031 -103 2065
rect -137 1963 -103 1997
rect -137 1895 -103 1929
rect -137 1827 -103 1861
rect -137 1759 -103 1793
rect -137 1691 -103 1725
rect -137 1623 -103 1657
rect -137 1555 -103 1589
rect -137 1487 -103 1521
rect -137 1419 -103 1453
rect -137 1351 -103 1385
rect -137 1283 -103 1317
rect -137 1215 -103 1249
rect -137 1147 -103 1181
rect -137 1079 -103 1113
rect -137 1011 -103 1045
rect -137 943 -103 977
rect -137 875 -103 909
rect -137 807 -103 841
rect -137 739 -103 773
rect -137 671 -103 705
rect -137 603 -103 637
rect -137 535 -103 569
rect -137 467 -103 501
rect -137 399 -103 433
rect -137 331 -103 365
rect -137 263 -103 297
rect -137 195 -103 229
rect -137 127 -103 161
rect -137 59 -103 93
rect -137 -9 -103 25
rect -137 -77 -103 -43
rect -137 -133 -103 -111
rect 6083 8974 6117 9003
rect 6083 8906 6117 8940
rect 6083 8838 6117 8872
rect 6083 8770 6117 8804
rect 6083 8702 6117 8736
rect 6083 8634 6117 8668
rect 6083 8566 6117 8600
rect 6083 8498 6117 8532
rect 6083 8430 6117 8464
rect 6083 8362 6117 8396
rect 6083 8294 6117 8328
rect 6083 8226 6117 8260
rect 6083 8158 6117 8192
rect 6083 8090 6117 8124
rect 6083 8022 6117 8056
rect 6083 7954 6117 7988
rect 6083 7886 6117 7920
rect 6083 7818 6117 7852
rect 6083 7750 6117 7784
rect 6083 7682 6117 7716
rect 6083 7614 6117 7648
rect 6083 7546 6117 7580
rect 6083 7478 6117 7512
rect 6083 7410 6117 7444
rect 6083 7342 6117 7376
rect 6083 7274 6117 7308
rect 6083 7206 6117 7240
rect 6083 7138 6117 7172
rect 6083 7070 6117 7104
rect 6083 7002 6117 7036
rect 6083 6934 6117 6968
rect 6083 6866 6117 6900
rect 6083 6798 6117 6832
rect 6083 6730 6117 6764
rect 6083 6662 6117 6696
rect 6083 6594 6117 6628
rect 6083 6526 6117 6560
rect 6083 6458 6117 6492
rect 6083 6390 6117 6424
rect 6083 6322 6117 6356
rect 6083 6254 6117 6288
rect 6083 6186 6117 6220
rect 6083 6118 6117 6152
rect 6083 6050 6117 6084
rect 6083 5982 6117 6016
rect 6083 5914 6117 5948
rect 6083 5846 6117 5880
rect 6083 5778 6117 5812
rect 6083 5710 6117 5744
rect 6083 5642 6117 5676
rect 6083 5574 6117 5608
rect 6083 5506 6117 5540
rect 6083 5438 6117 5472
rect 6083 5370 6117 5404
rect 6083 5302 6117 5336
rect 6083 5234 6117 5268
rect 6083 5166 6117 5200
rect 6083 5098 6117 5132
rect 6083 5030 6117 5064
rect 6083 4962 6117 4996
rect 6083 4894 6117 4928
rect 6083 4826 6117 4860
rect 6083 4758 6117 4792
rect 6083 4690 6117 4724
rect 6083 4622 6117 4656
rect 6083 4554 6117 4588
rect 6083 4486 6117 4520
rect 6083 4418 6117 4452
rect 6083 4350 6117 4384
rect 6083 4282 6117 4316
rect 6083 4214 6117 4248
rect 6083 4146 6117 4180
rect 6083 4078 6117 4112
rect 6083 4010 6117 4044
rect 6083 3942 6117 3976
rect 6083 3874 6117 3908
rect 6083 3806 6117 3840
rect 6083 3738 6117 3772
rect 6083 3670 6117 3704
rect 6083 3602 6117 3636
rect 6083 3534 6117 3568
rect 6083 3466 6117 3500
rect 6083 3398 6117 3432
rect 6083 3330 6117 3364
rect 6083 3262 6117 3296
rect 6083 3194 6117 3228
rect 6083 3126 6117 3160
rect 6083 3058 6117 3092
rect 6083 2990 6117 3024
rect 6083 2922 6117 2956
rect 6083 2854 6117 2888
rect 6083 2786 6117 2820
rect 6083 2718 6117 2752
rect 6083 2650 6117 2684
rect 6083 2582 6117 2616
rect 6083 2514 6117 2548
rect 6083 2446 6117 2480
rect 6083 2378 6117 2412
rect 6083 2310 6117 2344
rect 6083 2242 6117 2276
rect 6083 2174 6117 2208
rect 6083 2106 6117 2140
rect 6083 2038 6117 2072
rect 6083 1970 6117 2004
rect 6083 1902 6117 1936
rect 6083 1834 6117 1868
rect 6083 1766 6117 1800
rect 6083 1698 6117 1732
rect 6083 1630 6117 1664
rect 6083 1562 6117 1596
rect 6083 1494 6117 1528
rect 6083 1426 6117 1460
rect 6083 1358 6117 1392
rect 6083 1290 6117 1324
rect 6083 1222 6117 1256
rect 6083 1154 6117 1188
rect 6083 1086 6117 1120
rect 6083 1018 6117 1052
rect 6083 950 6117 984
rect 6083 882 6117 916
rect 6083 814 6117 848
rect 6083 746 6117 780
rect 6083 678 6117 712
rect 6083 610 6117 644
rect 6083 542 6117 576
rect 6083 474 6117 508
rect 6083 406 6117 440
rect 6083 338 6117 372
rect 6083 270 6117 304
rect 6083 202 6117 236
rect 6083 134 6117 168
rect 6083 66 6117 100
rect 6083 -2 6117 32
rect 6083 -70 6117 -36
rect 6083 -133 6117 -104
rect -137 -167 -33 -133
rect 1 -167 35 -133
rect 69 -167 103 -133
rect 137 -167 171 -133
rect 205 -167 239 -133
rect 273 -167 307 -133
rect 341 -167 375 -133
rect 409 -167 443 -133
rect 477 -167 511 -133
rect 545 -167 579 -133
rect 613 -167 647 -133
rect 681 -167 715 -133
rect 749 -167 783 -133
rect 817 -167 851 -133
rect 885 -167 919 -133
rect 953 -167 987 -133
rect 1021 -167 1055 -133
rect 1089 -167 1123 -133
rect 1157 -167 1191 -133
rect 1225 -167 1259 -133
rect 1293 -167 1327 -133
rect 1361 -167 1395 -133
rect 1429 -167 1463 -133
rect 1497 -167 1531 -133
rect 1565 -167 1599 -133
rect 1633 -167 1667 -133
rect 1701 -167 1735 -133
rect 1769 -167 1803 -133
rect 1837 -167 1871 -133
rect 1905 -167 1939 -133
rect 1973 -167 2007 -133
rect 2041 -167 2075 -133
rect 2109 -167 2143 -133
rect 2177 -167 2211 -133
rect 2245 -167 2279 -133
rect 2313 -167 2347 -133
rect 2381 -167 2415 -133
rect 2449 -167 2483 -133
rect 2517 -167 2551 -133
rect 2585 -167 2619 -133
rect 2653 -167 2687 -133
rect 2721 -167 2755 -133
rect 2789 -167 2823 -133
rect 2857 -167 2891 -133
rect 2925 -167 2959 -133
rect 2993 -167 3027 -133
rect 3061 -167 3095 -133
rect 3129 -167 3163 -133
rect 3197 -167 3231 -133
rect 3265 -167 3299 -133
rect 3333 -167 3367 -133
rect 3401 -167 3435 -133
rect 3469 -167 3503 -133
rect 3537 -167 3571 -133
rect 3605 -167 3639 -133
rect 3673 -167 3707 -133
rect 3741 -167 3775 -133
rect 3809 -167 3843 -133
rect 3877 -167 3911 -133
rect 3945 -167 3979 -133
rect 4013 -167 4047 -133
rect 4081 -167 4115 -133
rect 4149 -167 4183 -133
rect 4217 -167 4251 -133
rect 4285 -167 4319 -133
rect 4353 -167 4387 -133
rect 4421 -167 4455 -133
rect 4489 -167 4523 -133
rect 4557 -167 4591 -133
rect 4625 -167 4659 -133
rect 4693 -167 4727 -133
rect 4761 -167 4795 -133
rect 4829 -167 4863 -133
rect 4897 -167 4931 -133
rect 4965 -167 4999 -133
rect 5033 -167 5067 -133
rect 5101 -167 5135 -133
rect 5169 -167 5203 -133
rect 5237 -167 5271 -133
rect 5305 -167 5339 -133
rect 5373 -167 5407 -133
rect 5441 -167 5475 -133
rect 5509 -167 5543 -133
rect 5577 -167 5611 -133
rect 5645 -167 5679 -133
rect 5713 -167 5747 -133
rect 5781 -167 5815 -133
rect 5849 -167 5883 -133
rect 5917 -167 5951 -133
rect 5985 -167 6019 -133
rect 6053 -167 6117 -133
<< metal1 >>
rect 10 8850 90 9070
rect 310 8890 690 8970
rect 160 8846 240 8860
rect 310 8850 390 8890
rect 160 8794 174 8846
rect 226 8794 240 8846
rect 160 8766 240 8794
rect 160 8714 174 8766
rect 226 8714 240 8766
rect 160 8700 240 8714
rect 460 8846 540 8860
rect 610 8850 690 8890
rect 910 8890 1290 8970
rect 460 8794 474 8846
rect 526 8794 540 8846
rect 460 8766 540 8794
rect 460 8714 474 8766
rect 526 8714 540 8766
rect 460 8700 540 8714
rect 760 8846 840 8860
rect 910 8850 990 8890
rect 760 8794 774 8846
rect 826 8794 840 8846
rect 760 8766 840 8794
rect 760 8714 774 8766
rect 826 8714 840 8766
rect 760 8700 840 8714
rect 1060 8846 1140 8860
rect 1210 8850 1290 8890
rect 1510 8890 1890 8970
rect 1060 8794 1074 8846
rect 1126 8794 1140 8846
rect 1060 8766 1140 8794
rect 1060 8714 1074 8766
rect 1126 8714 1140 8766
rect 1060 8700 1140 8714
rect 1360 8846 1440 8860
rect 1510 8850 1590 8890
rect 1360 8794 1374 8846
rect 1426 8794 1440 8846
rect 1360 8766 1440 8794
rect 1360 8714 1374 8766
rect 1426 8714 1440 8766
rect 1360 8700 1440 8714
rect 1660 8846 1740 8860
rect 1810 8850 1890 8890
rect 2110 8890 2490 8970
rect 1660 8794 1674 8846
rect 1726 8794 1740 8846
rect 1660 8766 1740 8794
rect 1660 8714 1674 8766
rect 1726 8714 1740 8766
rect 1660 8700 1740 8714
rect 1960 8846 2040 8860
rect 2110 8850 2190 8890
rect 1960 8794 1974 8846
rect 2026 8794 2040 8846
rect 1960 8766 2040 8794
rect 1960 8714 1974 8766
rect 2026 8714 2040 8766
rect 1960 8700 2040 8714
rect 2260 8846 2340 8860
rect 2410 8850 2490 8890
rect 2710 8890 3090 8970
rect 2260 8794 2274 8846
rect 2326 8794 2340 8846
rect 2260 8766 2340 8794
rect 2260 8714 2274 8766
rect 2326 8714 2340 8766
rect 2260 8700 2340 8714
rect 2560 8846 2640 8860
rect 2710 8850 2790 8890
rect 2560 8794 2574 8846
rect 2626 8794 2640 8846
rect 2560 8766 2640 8794
rect 2560 8714 2574 8766
rect 2626 8714 2640 8766
rect 2560 8700 2640 8714
rect 2860 8846 2940 8860
rect 3010 8850 3090 8890
rect 3310 8890 3690 8970
rect 2860 8794 2874 8846
rect 2926 8794 2940 8846
rect 2860 8766 2940 8794
rect 2860 8714 2874 8766
rect 2926 8714 2940 8766
rect 2860 8700 2940 8714
rect 3160 8846 3240 8860
rect 3310 8850 3390 8890
rect 3160 8794 3174 8846
rect 3226 8794 3240 8846
rect 3160 8766 3240 8794
rect 3160 8714 3174 8766
rect 3226 8714 3240 8766
rect 3160 8700 3240 8714
rect 3460 8846 3540 8860
rect 3610 8850 3690 8890
rect 3910 8890 4290 8970
rect 3460 8794 3474 8846
rect 3526 8794 3540 8846
rect 3460 8766 3540 8794
rect 3460 8714 3474 8766
rect 3526 8714 3540 8766
rect 3460 8700 3540 8714
rect 3760 8846 3840 8860
rect 3910 8850 3990 8890
rect 3760 8794 3774 8846
rect 3826 8794 3840 8846
rect 3760 8766 3840 8794
rect 3760 8714 3774 8766
rect 3826 8714 3840 8766
rect 3760 8700 3840 8714
rect 4060 8846 4140 8860
rect 4210 8850 4290 8890
rect 4510 8890 4890 8970
rect 4060 8794 4074 8846
rect 4126 8794 4140 8846
rect 4060 8766 4140 8794
rect 4060 8714 4074 8766
rect 4126 8714 4140 8766
rect 4060 8700 4140 8714
rect 4360 8846 4440 8860
rect 4510 8850 4590 8890
rect 4360 8794 4374 8846
rect 4426 8794 4440 8846
rect 4360 8766 4440 8794
rect 4360 8714 4374 8766
rect 4426 8714 4440 8766
rect 4360 8700 4440 8714
rect 4660 8846 4740 8860
rect 4810 8850 4890 8890
rect 5110 8890 5490 8970
rect 4660 8794 4674 8846
rect 4726 8794 4740 8846
rect 4660 8766 4740 8794
rect 4660 8714 4674 8766
rect 4726 8714 4740 8766
rect 4660 8700 4740 8714
rect 4960 8846 5040 8860
rect 5110 8850 5190 8890
rect 4960 8794 4974 8846
rect 5026 8794 5040 8846
rect 4960 8766 5040 8794
rect 4960 8714 4974 8766
rect 5026 8714 5040 8766
rect 4960 8700 5040 8714
rect 5260 8846 5340 8860
rect 5410 8850 5490 8890
rect 5710 8890 5940 8970
rect 5260 8794 5274 8846
rect 5326 8794 5340 8846
rect 5260 8766 5340 8794
rect 5260 8714 5274 8766
rect 5326 8714 5340 8766
rect 5260 8700 5340 8714
rect 5560 8846 5640 8860
rect 5710 8850 5790 8890
rect 5560 8794 5574 8846
rect 5626 8794 5640 8846
rect 5860 8830 5940 8890
rect 5560 8766 5640 8794
rect 5560 8714 5574 8766
rect 5626 8714 5640 8766
rect 5560 8700 5640 8714
rect 160 146 240 160
rect 160 94 174 146
rect 226 94 240 146
rect 160 66 240 94
rect 10 -30 90 20
rect 160 14 174 66
rect 226 14 240 66
rect 160 0 240 14
rect 460 146 540 160
rect 460 94 474 146
rect 526 94 540 146
rect 460 66 540 94
rect 460 14 474 66
rect 526 14 540 66
rect 310 -30 390 10
rect 460 0 540 14
rect 760 146 840 160
rect 760 94 774 146
rect 826 94 840 146
rect 760 66 840 94
rect 760 14 774 66
rect 826 14 840 66
rect 10 -110 390 -30
rect 610 -30 690 10
rect 760 0 840 14
rect 1060 146 1140 160
rect 1060 94 1074 146
rect 1126 94 1140 146
rect 1060 66 1140 94
rect 1060 14 1074 66
rect 1126 14 1140 66
rect 910 -30 990 10
rect 1060 0 1140 14
rect 1360 146 1440 160
rect 1360 94 1374 146
rect 1426 94 1440 146
rect 1360 66 1440 94
rect 1360 14 1374 66
rect 1426 14 1440 66
rect 610 -110 990 -30
rect 1210 -30 1290 10
rect 1360 0 1440 14
rect 1660 146 1740 160
rect 1660 94 1674 146
rect 1726 94 1740 146
rect 1660 66 1740 94
rect 1660 14 1674 66
rect 1726 14 1740 66
rect 1510 -30 1590 10
rect 1660 0 1740 14
rect 1960 146 2040 160
rect 1960 94 1974 146
rect 2026 94 2040 146
rect 1960 66 2040 94
rect 1960 14 1974 66
rect 2026 14 2040 66
rect 1210 -110 1590 -30
rect 1810 -30 1890 10
rect 1960 0 2040 14
rect 2260 146 2340 160
rect 2260 94 2274 146
rect 2326 94 2340 146
rect 2260 66 2340 94
rect 2260 14 2274 66
rect 2326 14 2340 66
rect 2110 -30 2190 10
rect 2260 0 2340 14
rect 2560 146 2640 160
rect 2560 94 2574 146
rect 2626 94 2640 146
rect 2560 66 2640 94
rect 2560 14 2574 66
rect 2626 14 2640 66
rect 1810 -110 2190 -30
rect 2410 -30 2490 10
rect 2560 0 2640 14
rect 2860 146 2940 160
rect 2860 94 2874 146
rect 2926 94 2940 146
rect 2860 66 2940 94
rect 2860 14 2874 66
rect 2926 14 2940 66
rect 2710 -30 2790 10
rect 2860 0 2940 14
rect 3160 146 3240 160
rect 3160 94 3174 146
rect 3226 94 3240 146
rect 3160 66 3240 94
rect 3160 14 3174 66
rect 3226 14 3240 66
rect 2410 -110 2790 -30
rect 3010 -30 3090 10
rect 3160 0 3240 14
rect 3460 146 3540 160
rect 3460 94 3474 146
rect 3526 94 3540 146
rect 3460 66 3540 94
rect 3460 14 3474 66
rect 3526 14 3540 66
rect 3310 -30 3390 10
rect 3460 0 3540 14
rect 3760 146 3840 160
rect 3760 94 3774 146
rect 3826 94 3840 146
rect 3760 66 3840 94
rect 3760 14 3774 66
rect 3826 14 3840 66
rect 3010 -110 3390 -30
rect 3610 -30 3690 10
rect 3760 0 3840 14
rect 4060 146 4140 160
rect 4060 94 4074 146
rect 4126 94 4140 146
rect 4060 66 4140 94
rect 4060 14 4074 66
rect 4126 14 4140 66
rect 3910 -30 3990 10
rect 4060 0 4140 14
rect 4360 146 4440 160
rect 4360 94 4374 146
rect 4426 94 4440 146
rect 4360 66 4440 94
rect 4360 14 4374 66
rect 4426 14 4440 66
rect 3610 -110 3990 -30
rect 4210 -30 4290 10
rect 4360 0 4440 14
rect 4660 146 4740 160
rect 4660 94 4674 146
rect 4726 94 4740 146
rect 4660 66 4740 94
rect 4660 14 4674 66
rect 4726 14 4740 66
rect 4510 -30 4590 10
rect 4660 0 4740 14
rect 4960 146 5040 160
rect 4960 94 4974 146
rect 5026 94 5040 146
rect 4960 66 5040 94
rect 4960 14 4974 66
rect 5026 14 5040 66
rect 4210 -110 4590 -30
rect 4810 -30 4890 10
rect 4960 0 5040 14
rect 5260 146 5340 160
rect 5260 94 5274 146
rect 5326 94 5340 146
rect 5260 66 5340 94
rect 5260 14 5274 66
rect 5326 14 5340 66
rect 5110 -30 5190 10
rect 5260 0 5340 14
rect 5560 146 5640 160
rect 5560 94 5574 146
rect 5626 94 5640 146
rect 5560 66 5640 94
rect 5560 14 5574 66
rect 5626 14 5640 66
rect 4810 -110 5190 -30
rect 5410 -30 5490 10
rect 5560 0 5640 14
rect 5860 146 5940 160
rect 5860 94 5874 146
rect 5926 94 5940 146
rect 5860 66 5940 94
rect 5860 14 5874 66
rect 5926 14 5940 66
rect 5710 -30 5790 10
rect 5860 0 5940 14
rect 5410 -110 5790 -30
<< via1 >>
rect 174 8794 226 8846
rect 174 8714 226 8766
rect 474 8794 526 8846
rect 474 8714 526 8766
rect 774 8794 826 8846
rect 774 8714 826 8766
rect 1074 8794 1126 8846
rect 1074 8714 1126 8766
rect 1374 8794 1426 8846
rect 1374 8714 1426 8766
rect 1674 8794 1726 8846
rect 1674 8714 1726 8766
rect 1974 8794 2026 8846
rect 1974 8714 2026 8766
rect 2274 8794 2326 8846
rect 2274 8714 2326 8766
rect 2574 8794 2626 8846
rect 2574 8714 2626 8766
rect 2874 8794 2926 8846
rect 2874 8714 2926 8766
rect 3174 8794 3226 8846
rect 3174 8714 3226 8766
rect 3474 8794 3526 8846
rect 3474 8714 3526 8766
rect 3774 8794 3826 8846
rect 3774 8714 3826 8766
rect 4074 8794 4126 8846
rect 4074 8714 4126 8766
rect 4374 8794 4426 8846
rect 4374 8714 4426 8766
rect 4674 8794 4726 8846
rect 4674 8714 4726 8766
rect 4974 8794 5026 8846
rect 4974 8714 5026 8766
rect 5274 8794 5326 8846
rect 5274 8714 5326 8766
rect 5574 8794 5626 8846
rect 5574 8714 5626 8766
rect 174 94 226 146
rect 174 14 226 66
rect 474 94 526 146
rect 474 14 526 66
rect 774 94 826 146
rect 774 14 826 66
rect 1074 94 1126 146
rect 1074 14 1126 66
rect 1374 94 1426 146
rect 1374 14 1426 66
rect 1674 94 1726 146
rect 1674 14 1726 66
rect 1974 94 2026 146
rect 1974 14 2026 66
rect 2274 94 2326 146
rect 2274 14 2326 66
rect 2574 94 2626 146
rect 2574 14 2626 66
rect 2874 94 2926 146
rect 2874 14 2926 66
rect 3174 94 3226 146
rect 3174 14 3226 66
rect 3474 94 3526 146
rect 3474 14 3526 66
rect 3774 94 3826 146
rect 3774 14 3826 66
rect 4074 94 4126 146
rect 4074 14 4126 66
rect 4374 94 4426 146
rect 4374 14 4426 66
rect 4674 94 4726 146
rect 4674 14 4726 66
rect 4974 94 5026 146
rect 4974 14 5026 66
rect 5274 94 5326 146
rect 5274 14 5326 66
rect 5574 94 5626 146
rect 5574 14 5626 66
rect 5874 94 5926 146
rect 5874 14 5926 66
<< metal2 >>
rect 160 8846 240 9070
rect 160 8794 174 8846
rect 226 8794 240 8846
rect 160 8766 240 8794
rect 160 8714 174 8766
rect 226 8714 240 8766
rect 160 8700 240 8714
rect 460 8890 840 8970
rect 460 8846 540 8890
rect 460 8794 474 8846
rect 526 8794 540 8846
rect 460 8766 540 8794
rect 460 8714 474 8766
rect 526 8714 540 8766
rect 460 8700 540 8714
rect 760 8846 840 8890
rect 760 8794 774 8846
rect 826 8794 840 8846
rect 760 8766 840 8794
rect 760 8714 774 8766
rect 826 8714 840 8766
rect 760 8700 840 8714
rect 1060 8890 1440 8970
rect 1060 8846 1140 8890
rect 1060 8794 1074 8846
rect 1126 8794 1140 8846
rect 1060 8766 1140 8794
rect 1060 8714 1074 8766
rect 1126 8714 1140 8766
rect 1060 8700 1140 8714
rect 1360 8846 1440 8890
rect 1360 8794 1374 8846
rect 1426 8794 1440 8846
rect 1360 8766 1440 8794
rect 1360 8714 1374 8766
rect 1426 8714 1440 8766
rect 1360 8700 1440 8714
rect 1660 8890 2040 8970
rect 1660 8846 1740 8890
rect 1660 8794 1674 8846
rect 1726 8794 1740 8846
rect 1660 8766 1740 8794
rect 1660 8714 1674 8766
rect 1726 8714 1740 8766
rect 1660 8700 1740 8714
rect 1960 8846 2040 8890
rect 1960 8794 1974 8846
rect 2026 8794 2040 8846
rect 1960 8766 2040 8794
rect 1960 8714 1974 8766
rect 2026 8714 2040 8766
rect 1960 8700 2040 8714
rect 2260 8890 2640 8970
rect 2260 8846 2340 8890
rect 2260 8794 2274 8846
rect 2326 8794 2340 8846
rect 2260 8766 2340 8794
rect 2260 8714 2274 8766
rect 2326 8714 2340 8766
rect 2260 8700 2340 8714
rect 2560 8846 2640 8890
rect 2560 8794 2574 8846
rect 2626 8794 2640 8846
rect 2560 8766 2640 8794
rect 2560 8714 2574 8766
rect 2626 8714 2640 8766
rect 2560 8700 2640 8714
rect 2860 8890 3240 8970
rect 2860 8846 2940 8890
rect 2860 8794 2874 8846
rect 2926 8794 2940 8846
rect 2860 8766 2940 8794
rect 2860 8714 2874 8766
rect 2926 8714 2940 8766
rect 2860 8700 2940 8714
rect 3160 8846 3240 8890
rect 3160 8794 3174 8846
rect 3226 8794 3240 8846
rect 3160 8766 3240 8794
rect 3160 8714 3174 8766
rect 3226 8714 3240 8766
rect 3160 8700 3240 8714
rect 3460 8890 3840 8970
rect 3460 8846 3540 8890
rect 3460 8794 3474 8846
rect 3526 8794 3540 8846
rect 3460 8766 3540 8794
rect 3460 8714 3474 8766
rect 3526 8714 3540 8766
rect 3460 8700 3540 8714
rect 3760 8846 3840 8890
rect 3760 8794 3774 8846
rect 3826 8794 3840 8846
rect 3760 8766 3840 8794
rect 3760 8714 3774 8766
rect 3826 8714 3840 8766
rect 3760 8700 3840 8714
rect 4060 8890 4440 8970
rect 4060 8846 4140 8890
rect 4060 8794 4074 8846
rect 4126 8794 4140 8846
rect 4060 8766 4140 8794
rect 4060 8714 4074 8766
rect 4126 8714 4140 8766
rect 4060 8700 4140 8714
rect 4360 8846 4440 8890
rect 4360 8794 4374 8846
rect 4426 8794 4440 8846
rect 4360 8766 4440 8794
rect 4360 8714 4374 8766
rect 4426 8714 4440 8766
rect 4360 8700 4440 8714
rect 4660 8890 5040 8970
rect 4660 8846 4740 8890
rect 4660 8794 4674 8846
rect 4726 8794 4740 8846
rect 4660 8766 4740 8794
rect 4660 8714 4674 8766
rect 4726 8714 4740 8766
rect 4660 8700 4740 8714
rect 4960 8846 5040 8890
rect 4960 8794 4974 8846
rect 5026 8794 5040 8846
rect 4960 8766 5040 8794
rect 4960 8714 4974 8766
rect 5026 8714 5040 8766
rect 4960 8700 5040 8714
rect 5260 8890 5640 8970
rect 5260 8846 5340 8890
rect 5260 8794 5274 8846
rect 5326 8794 5340 8846
rect 5260 8766 5340 8794
rect 5260 8714 5274 8766
rect 5326 8714 5340 8766
rect 5260 8700 5340 8714
rect 5560 8846 5640 8890
rect 5560 8794 5574 8846
rect 5626 8794 5640 8846
rect 5560 8766 5640 8794
rect 5560 8714 5574 8766
rect 5626 8714 5640 8766
rect 5560 8700 5640 8714
rect 160 146 240 160
rect 160 94 174 146
rect 226 94 240 146
rect 160 66 240 94
rect 160 14 174 66
rect 226 14 240 66
rect 160 -30 240 14
rect 460 146 540 160
rect 460 94 474 146
rect 526 94 540 146
rect 460 66 540 94
rect 460 14 474 66
rect 526 14 540 66
rect 460 -30 540 14
rect 160 -110 540 -30
rect 760 146 840 160
rect 760 94 774 146
rect 826 94 840 146
rect 760 66 840 94
rect 760 14 774 66
rect 826 14 840 66
rect 760 -30 840 14
rect 1060 146 1140 160
rect 1060 94 1074 146
rect 1126 94 1140 146
rect 1060 66 1140 94
rect 1060 14 1074 66
rect 1126 14 1140 66
rect 1060 -30 1140 14
rect 760 -110 1140 -30
rect 1360 146 1440 160
rect 1360 94 1374 146
rect 1426 94 1440 146
rect 1360 66 1440 94
rect 1360 14 1374 66
rect 1426 14 1440 66
rect 1360 -30 1440 14
rect 1660 146 1740 160
rect 1660 94 1674 146
rect 1726 94 1740 146
rect 1660 66 1740 94
rect 1660 14 1674 66
rect 1726 14 1740 66
rect 1660 -30 1740 14
rect 1360 -110 1740 -30
rect 1960 146 2040 160
rect 1960 94 1974 146
rect 2026 94 2040 146
rect 1960 66 2040 94
rect 1960 14 1974 66
rect 2026 14 2040 66
rect 1960 -30 2040 14
rect 2260 146 2340 160
rect 2260 94 2274 146
rect 2326 94 2340 146
rect 2260 66 2340 94
rect 2260 14 2274 66
rect 2326 14 2340 66
rect 2260 -30 2340 14
rect 1960 -110 2340 -30
rect 2560 146 2640 160
rect 2560 94 2574 146
rect 2626 94 2640 146
rect 2560 66 2640 94
rect 2560 14 2574 66
rect 2626 14 2640 66
rect 2560 -30 2640 14
rect 2860 146 2940 160
rect 2860 94 2874 146
rect 2926 94 2940 146
rect 2860 66 2940 94
rect 2860 14 2874 66
rect 2926 14 2940 66
rect 2860 -30 2940 14
rect 2560 -110 2940 -30
rect 3160 146 3240 160
rect 3160 94 3174 146
rect 3226 94 3240 146
rect 3160 66 3240 94
rect 3160 14 3174 66
rect 3226 14 3240 66
rect 3160 -30 3240 14
rect 3460 146 3540 160
rect 3460 94 3474 146
rect 3526 94 3540 146
rect 3460 66 3540 94
rect 3460 14 3474 66
rect 3526 14 3540 66
rect 3460 -30 3540 14
rect 3160 -110 3540 -30
rect 3760 146 3840 160
rect 3760 94 3774 146
rect 3826 94 3840 146
rect 3760 66 3840 94
rect 3760 14 3774 66
rect 3826 14 3840 66
rect 3760 -30 3840 14
rect 4060 146 4140 160
rect 4060 94 4074 146
rect 4126 94 4140 146
rect 4060 66 4140 94
rect 4060 14 4074 66
rect 4126 14 4140 66
rect 4060 -30 4140 14
rect 3760 -110 4140 -30
rect 4360 146 4440 160
rect 4360 94 4374 146
rect 4426 94 4440 146
rect 4360 66 4440 94
rect 4360 14 4374 66
rect 4426 14 4440 66
rect 4360 -30 4440 14
rect 4660 146 4740 160
rect 4660 94 4674 146
rect 4726 94 4740 146
rect 4660 66 4740 94
rect 4660 14 4674 66
rect 4726 14 4740 66
rect 4660 -30 4740 14
rect 4360 -110 4740 -30
rect 4960 146 5040 160
rect 4960 94 4974 146
rect 5026 94 5040 146
rect 4960 66 5040 94
rect 4960 14 4974 66
rect 5026 14 5040 66
rect 4960 -30 5040 14
rect 5260 146 5340 160
rect 5260 94 5274 146
rect 5326 94 5340 146
rect 5260 66 5340 94
rect 5260 14 5274 66
rect 5326 14 5340 66
rect 5260 -30 5340 14
rect 4960 -110 5340 -30
rect 5560 146 5640 160
rect 5560 94 5574 146
rect 5626 94 5640 146
rect 5560 66 5640 94
rect 5560 14 5574 66
rect 5626 14 5640 66
rect 5560 -30 5640 14
rect 5860 146 5940 160
rect 5860 94 5874 146
rect 5926 94 5940 146
rect 5860 66 5940 94
rect 5860 14 5874 66
rect 5926 14 5940 66
rect 5860 -30 5940 14
rect 5560 -110 5940 -30
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_0
timestamp 1757161594
transform 1 0 2300 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_1
timestamp 1757161594
transform 1 0 1850 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_2
timestamp 1757161594
transform 1 0 2000 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_3
timestamp 1757161594
transform 1 0 2150 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_4
timestamp 1757161594
transform 1 0 1700 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_5
timestamp 1757161594
transform 1 0 1550 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_6
timestamp 1757161594
transform 1 0 1400 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_7
timestamp 1757161594
transform 1 0 1250 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_8
timestamp 1757161594
transform 1 0 650 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_9
timestamp 1757161594
transform 1 0 800 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_10
timestamp 1757161594
transform 1 0 950 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_11
timestamp 1757161594
transform 1 0 1100 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_12
timestamp 1757161594
transform 1 0 500 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_13
timestamp 1757161594
transform 1 0 350 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_14
timestamp 1757161594
transform 1 0 200 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_15
timestamp 1757161594
transform 1 0 50 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_16
timestamp 1757161594
transform 1 0 3650 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_17
timestamp 1757161594
transform 1 0 3800 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_18
timestamp 1757161594
transform 1 0 3950 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_19
timestamp 1757161594
transform 1 0 4100 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_20
timestamp 1757161594
transform 1 0 4250 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_21
timestamp 1757161594
transform 1 0 4400 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_22
timestamp 1757161594
transform 1 0 4550 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_23
timestamp 1757161594
transform 1 0 4700 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_24
timestamp 1757161594
transform 1 0 2450 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_25
timestamp 1757161594
transform 1 0 2600 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_26
timestamp 1757161594
transform 1 0 2750 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_27
timestamp 1757161594
transform 1 0 2900 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_28
timestamp 1757161594
transform 1 0 3050 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_29
timestamp 1757161594
transform 1 0 3200 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_30
timestamp 1757161594
transform 1 0 3350 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_31
timestamp 1757161594
transform 1 0 3500 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_32
timestamp 1757161594
transform 1 0 4850 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_33
timestamp 1757161594
transform 1 0 5000 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_34
timestamp 1757161594
transform 1 0 5150 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_35
timestamp 1757161594
transform 1 0 5300 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_36
timestamp 1757161594
transform 1 0 5450 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_37
timestamp 1757161594
transform 1 0 5600 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_38
timestamp 1757161594
transform 1 0 5750 0 1 4430
box -50 -4430 50 4430
use sky130_fd_pr__res_generic_po_RETGBZ  sky130_fd_pr__res_generic_po_RETGBZ_40
timestamp 1757161594
transform 1 0 5900 0 1 4430
box -50 -4430 50 4430
<< end >>
