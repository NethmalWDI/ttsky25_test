magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -184 -117 184 55
<< nmoslvt >>
rect -100 -91 100 29
<< ndiff >>
rect -158 -14 -100 29
rect -158 -48 -146 -14
rect -112 -48 -100 -14
rect -158 -91 -100 -48
rect 100 -14 158 29
rect 100 -48 112 -14
rect 146 -48 158 -14
rect 100 -91 158 -48
<< ndiffc >>
rect -146 -48 -112 -14
rect 112 -48 146 -14
<< poly >>
rect -75 101 75 117
rect -75 84 -51 101
rect -100 67 -51 84
rect -17 67 17 101
rect 51 84 75 101
rect 51 67 100 84
rect -100 29 100 67
rect -100 -117 100 -91
<< polycont >>
rect -51 67 -17 101
rect 17 67 51 101
<< locali >>
rect -75 67 -53 101
rect -17 67 17 101
rect 53 67 75 101
rect -146 -14 -112 19
rect -146 -81 -112 -48
rect 112 -14 146 19
rect 112 -81 146 -48
<< viali >>
rect -53 67 -51 101
rect -51 67 -19 101
rect 19 67 51 101
rect 51 67 53 101
rect -146 -48 -112 -14
rect 112 -48 146 -14
<< metal1 >>
rect -71 101 71 107
rect -71 67 -53 101
rect -19 67 19 101
rect 53 67 71 101
rect -71 61 71 67
rect -152 -14 -106 15
rect -152 -48 -146 -14
rect -112 -48 -106 -14
rect -152 -77 -106 -48
rect 106 -14 152 15
rect 106 -48 112 -14
rect 146 -48 152 -14
rect 106 -77 152 -48
<< end >>
