magic
tech sky130A
magscale 1 2
timestamp 1757161594
<< pwell >>
rect -1084 -257 1084 195
<< nmoslvt >>
rect -1000 -231 1000 169
<< ndiff >>
rect -1058 88 -1000 169
rect -1058 54 -1046 88
rect -1012 54 -1000 88
rect -1058 20 -1000 54
rect -1058 -14 -1046 20
rect -1012 -14 -1000 20
rect -1058 -48 -1000 -14
rect -1058 -82 -1046 -48
rect -1012 -82 -1000 -48
rect -1058 -116 -1000 -82
rect -1058 -150 -1046 -116
rect -1012 -150 -1000 -116
rect -1058 -231 -1000 -150
rect 1000 88 1058 169
rect 1000 54 1012 88
rect 1046 54 1058 88
rect 1000 20 1058 54
rect 1000 -14 1012 20
rect 1046 -14 1058 20
rect 1000 -48 1058 -14
rect 1000 -82 1012 -48
rect 1046 -82 1058 -48
rect 1000 -116 1058 -82
rect 1000 -150 1012 -116
rect 1046 -150 1058 -116
rect 1000 -231 1058 -150
<< ndiffc >>
rect -1046 54 -1012 88
rect -1046 -14 -1012 20
rect -1046 -82 -1012 -48
rect -1046 -150 -1012 -116
rect 1012 54 1046 88
rect 1012 -14 1046 20
rect 1012 -82 1046 -48
rect 1012 -150 1046 -116
<< poly >>
rect -705 241 705 257
rect -705 224 -663 241
rect -1000 207 -663 224
rect -629 207 -595 241
rect -561 207 -527 241
rect -493 207 -459 241
rect -425 207 -391 241
rect -357 207 -323 241
rect -289 207 -255 241
rect -221 207 -187 241
rect -153 207 -119 241
rect -85 207 -51 241
rect -17 207 17 241
rect 51 207 85 241
rect 119 207 153 241
rect 187 207 221 241
rect 255 207 289 241
rect 323 207 357 241
rect 391 207 425 241
rect 459 207 493 241
rect 527 207 561 241
rect 595 207 629 241
rect 663 224 705 241
rect 663 207 1000 224
rect -1000 169 1000 207
rect -1000 -257 1000 -231
<< polycont >>
rect -663 207 -629 241
rect -595 207 -561 241
rect -527 207 -493 241
rect -459 207 -425 241
rect -391 207 -357 241
rect -323 207 -289 241
rect -255 207 -221 241
rect -187 207 -153 241
rect -119 207 -85 241
rect -51 207 -17 241
rect 17 207 51 241
rect 85 207 119 241
rect 153 207 187 241
rect 221 207 255 241
rect 289 207 323 241
rect 357 207 391 241
rect 425 207 459 241
rect 493 207 527 241
rect 561 207 595 241
rect 629 207 663 241
<< locali >>
rect -705 207 -665 241
rect -629 207 -595 241
rect -559 207 -527 241
rect -487 207 -459 241
rect -415 207 -391 241
rect -343 207 -323 241
rect -271 207 -255 241
rect -199 207 -187 241
rect -127 207 -119 241
rect -55 207 -51 241
rect 51 207 55 241
rect 119 207 127 241
rect 187 207 199 241
rect 255 207 271 241
rect 323 207 343 241
rect 391 207 415 241
rect 459 207 487 241
rect 527 207 559 241
rect 595 207 629 241
rect 665 207 705 241
rect -1046 94 -1012 117
rect -1046 22 -1012 54
rect -1046 -48 -1012 -14
rect -1046 -116 -1012 -84
rect -1046 -179 -1012 -156
rect 1012 94 1046 117
rect 1012 22 1046 54
rect 1012 -48 1046 -14
rect 1012 -116 1046 -84
rect 1012 -179 1046 -156
<< viali >>
rect -665 207 -663 241
rect -663 207 -631 241
rect -593 207 -561 241
rect -561 207 -559 241
rect -521 207 -493 241
rect -493 207 -487 241
rect -449 207 -425 241
rect -425 207 -415 241
rect -377 207 -357 241
rect -357 207 -343 241
rect -305 207 -289 241
rect -289 207 -271 241
rect -233 207 -221 241
rect -221 207 -199 241
rect -161 207 -153 241
rect -153 207 -127 241
rect -89 207 -85 241
rect -85 207 -55 241
rect -17 207 17 241
rect 55 207 85 241
rect 85 207 89 241
rect 127 207 153 241
rect 153 207 161 241
rect 199 207 221 241
rect 221 207 233 241
rect 271 207 289 241
rect 289 207 305 241
rect 343 207 357 241
rect 357 207 377 241
rect 415 207 425 241
rect 425 207 449 241
rect 487 207 493 241
rect 493 207 521 241
rect 559 207 561 241
rect 561 207 593 241
rect 631 207 663 241
rect 663 207 665 241
rect -1046 88 -1012 94
rect -1046 60 -1012 88
rect -1046 20 -1012 22
rect -1046 -12 -1012 20
rect -1046 -82 -1012 -50
rect -1046 -84 -1012 -82
rect -1046 -150 -1012 -122
rect -1046 -156 -1012 -150
rect 1012 88 1046 94
rect 1012 60 1046 88
rect 1012 20 1046 22
rect 1012 -12 1046 20
rect 1012 -82 1046 -50
rect 1012 -84 1046 -82
rect 1012 -150 1046 -122
rect 1012 -156 1046 -150
<< metal1 >>
rect -701 241 701 247
rect -701 207 -665 241
rect -631 207 -593 241
rect -559 207 -521 241
rect -487 207 -449 241
rect -415 207 -377 241
rect -343 207 -305 241
rect -271 207 -233 241
rect -199 207 -161 241
rect -127 207 -89 241
rect -55 207 -17 241
rect 17 207 55 241
rect 89 207 127 241
rect 161 207 199 241
rect 233 207 271 241
rect 305 207 343 241
rect 377 207 415 241
rect 449 207 487 241
rect 521 207 559 241
rect 593 207 631 241
rect 665 207 701 241
rect -701 201 701 207
rect -1052 94 -1006 113
rect -1052 60 -1046 94
rect -1012 60 -1006 94
rect -1052 22 -1006 60
rect -1052 -12 -1046 22
rect -1012 -12 -1006 22
rect -1052 -50 -1006 -12
rect -1052 -84 -1046 -50
rect -1012 -84 -1006 -50
rect -1052 -122 -1006 -84
rect -1052 -156 -1046 -122
rect -1012 -156 -1006 -122
rect -1052 -175 -1006 -156
rect 1006 94 1052 113
rect 1006 60 1012 94
rect 1046 60 1052 94
rect 1006 22 1052 60
rect 1006 -12 1012 22
rect 1046 -12 1052 22
rect 1006 -50 1052 -12
rect 1006 -84 1012 -50
rect 1046 -84 1052 -50
rect 1006 -122 1052 -84
rect 1006 -156 1012 -122
rect 1046 -156 1052 -122
rect 1006 -175 1052 -156
<< end >>
